module PositDivSqrter15_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [14:0] io_A,
  input  [14:0] io_B,
  output        io_diviValid,
  output        io_sqrtValid,
  output        io_invalidExc,
  output [14:0] io_Q
);
  reg [3:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [6:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [10:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [14:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [14:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [12:0] _T_4; // @[convert.scala 19:24]
  wire [12:0] _T_5; // @[convert.scala 19:43]
  wire [12:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [4:0] _T_68; // @[LZD.scala 44:32]
  wire [3:0] _T_69; // @[LZD.scala 43:32]
  wire [1:0] _T_70; // @[LZD.scala 43:32]
  wire  _T_71; // @[LZD.scala 39:14]
  wire  _T_72; // @[LZD.scala 39:21]
  wire  _T_73; // @[LZD.scala 39:30]
  wire  _T_74; // @[LZD.scala 39:27]
  wire  _T_75; // @[LZD.scala 39:25]
  wire [1:0] _T_76; // @[Cat.scala 29:58]
  wire [1:0] _T_77; // @[LZD.scala 44:32]
  wire  _T_78; // @[LZD.scala 39:14]
  wire  _T_79; // @[LZD.scala 39:21]
  wire  _T_80; // @[LZD.scala 39:30]
  wire  _T_81; // @[LZD.scala 39:27]
  wire  _T_82; // @[LZD.scala 39:25]
  wire [1:0] _T_83; // @[Cat.scala 29:58]
  wire  _T_84; // @[Shift.scala 12:21]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[LZD.scala 49:16]
  wire  _T_87; // @[LZD.scala 49:27]
  wire  _T_88; // @[LZD.scala 49:25]
  wire  _T_89; // @[LZD.scala 49:47]
  wire  _T_90; // @[LZD.scala 49:59]
  wire  _T_91; // @[LZD.scala 49:35]
  wire [2:0] _T_93; // @[Cat.scala 29:58]
  wire  _T_94; // @[LZD.scala 44:32]
  wire  _T_96; // @[Shift.scala 12:21]
  wire [1:0] _T_98; // @[Cat.scala 29:58]
  wire [1:0] _T_99; // @[LZD.scala 55:32]
  wire [1:0] _T_100; // @[LZD.scala 55:20]
  wire [2:0] _T_101; // @[Cat.scala 29:58]
  wire  _T_102; // @[Shift.scala 12:21]
  wire [2:0] _T_104; // @[LZD.scala 55:32]
  wire [2:0] _T_105; // @[LZD.scala 55:20]
  wire [3:0] _T_106; // @[Cat.scala 29:58]
  wire [3:0] _T_107; // @[convert.scala 21:22]
  wire [11:0] _T_108; // @[convert.scala 22:36]
  wire  _T_109; // @[Shift.scala 16:24]
  wire  _T_111; // @[Shift.scala 12:21]
  wire [3:0] _T_112; // @[Shift.scala 64:52]
  wire [11:0] _T_114; // @[Cat.scala 29:58]
  wire [11:0] _T_115; // @[Shift.scala 64:27]
  wire [2:0] _T_116; // @[Shift.scala 66:70]
  wire  _T_117; // @[Shift.scala 12:21]
  wire [7:0] _T_118; // @[Shift.scala 64:52]
  wire [11:0] _T_120; // @[Cat.scala 29:58]
  wire [11:0] _T_121; // @[Shift.scala 64:27]
  wire [1:0] _T_122; // @[Shift.scala 66:70]
  wire  _T_123; // @[Shift.scala 12:21]
  wire [9:0] _T_124; // @[Shift.scala 64:52]
  wire [11:0] _T_126; // @[Cat.scala 29:58]
  wire [11:0] _T_127; // @[Shift.scala 64:27]
  wire  _T_128; // @[Shift.scala 66:70]
  wire [10:0] _T_130; // @[Shift.scala 64:52]
  wire [11:0] _T_131; // @[Cat.scala 29:58]
  wire [11:0] _T_132; // @[Shift.scala 64:27]
  wire [11:0] _T_133; // @[Shift.scala 16:10]
  wire  _T_134; // @[convert.scala 23:34]
  wire [10:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_136; // @[convert.scala 25:26]
  wire [3:0] _T_138; // @[convert.scala 25:42]
  wire  _T_141; // @[convert.scala 26:67]
  wire  _T_142; // @[convert.scala 26:51]
  wire [5:0] _T_143; // @[Cat.scala 29:58]
  wire [13:0] _T_145; // @[convert.scala 29:56]
  wire  _T_146; // @[convert.scala 29:60]
  wire  _T_147; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_150; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_159; // @[convert.scala 18:24]
  wire  _T_160; // @[convert.scala 18:40]
  wire  _T_161; // @[convert.scala 18:36]
  wire [12:0] _T_162; // @[convert.scala 19:24]
  wire [12:0] _T_163; // @[convert.scala 19:43]
  wire [12:0] _T_164; // @[convert.scala 19:39]
  wire [7:0] _T_165; // @[LZD.scala 43:32]
  wire [3:0] _T_166; // @[LZD.scala 43:32]
  wire [1:0] _T_167; // @[LZD.scala 43:32]
  wire  _T_168; // @[LZD.scala 39:14]
  wire  _T_169; // @[LZD.scala 39:21]
  wire  _T_170; // @[LZD.scala 39:30]
  wire  _T_171; // @[LZD.scala 39:27]
  wire  _T_172; // @[LZD.scala 39:25]
  wire [1:0] _T_173; // @[Cat.scala 29:58]
  wire [1:0] _T_174; // @[LZD.scala 44:32]
  wire  _T_175; // @[LZD.scala 39:14]
  wire  _T_176; // @[LZD.scala 39:21]
  wire  _T_177; // @[LZD.scala 39:30]
  wire  _T_178; // @[LZD.scala 39:27]
  wire  _T_179; // @[LZD.scala 39:25]
  wire [1:0] _T_180; // @[Cat.scala 29:58]
  wire  _T_181; // @[Shift.scala 12:21]
  wire  _T_182; // @[Shift.scala 12:21]
  wire  _T_183; // @[LZD.scala 49:16]
  wire  _T_184; // @[LZD.scala 49:27]
  wire  _T_185; // @[LZD.scala 49:25]
  wire  _T_186; // @[LZD.scala 49:47]
  wire  _T_187; // @[LZD.scala 49:59]
  wire  _T_188; // @[LZD.scala 49:35]
  wire [2:0] _T_190; // @[Cat.scala 29:58]
  wire [3:0] _T_191; // @[LZD.scala 44:32]
  wire [1:0] _T_192; // @[LZD.scala 43:32]
  wire  _T_193; // @[LZD.scala 39:14]
  wire  _T_194; // @[LZD.scala 39:21]
  wire  _T_195; // @[LZD.scala 39:30]
  wire  _T_196; // @[LZD.scala 39:27]
  wire  _T_197; // @[LZD.scala 39:25]
  wire [1:0] _T_198; // @[Cat.scala 29:58]
  wire [1:0] _T_199; // @[LZD.scala 44:32]
  wire  _T_200; // @[LZD.scala 39:14]
  wire  _T_201; // @[LZD.scala 39:21]
  wire  _T_202; // @[LZD.scala 39:30]
  wire  _T_203; // @[LZD.scala 39:27]
  wire  _T_204; // @[LZD.scala 39:25]
  wire [1:0] _T_205; // @[Cat.scala 29:58]
  wire  _T_206; // @[Shift.scala 12:21]
  wire  _T_207; // @[Shift.scala 12:21]
  wire  _T_208; // @[LZD.scala 49:16]
  wire  _T_209; // @[LZD.scala 49:27]
  wire  _T_210; // @[LZD.scala 49:25]
  wire  _T_211; // @[LZD.scala 49:47]
  wire  _T_212; // @[LZD.scala 49:59]
  wire  _T_213; // @[LZD.scala 49:35]
  wire [2:0] _T_215; // @[Cat.scala 29:58]
  wire  _T_216; // @[Shift.scala 12:21]
  wire  _T_217; // @[Shift.scala 12:21]
  wire  _T_218; // @[LZD.scala 49:16]
  wire  _T_219; // @[LZD.scala 49:27]
  wire  _T_220; // @[LZD.scala 49:25]
  wire [1:0] _T_221; // @[LZD.scala 49:47]
  wire [1:0] _T_222; // @[LZD.scala 49:59]
  wire [1:0] _T_223; // @[LZD.scala 49:35]
  wire [3:0] _T_225; // @[Cat.scala 29:58]
  wire [4:0] _T_226; // @[LZD.scala 44:32]
  wire [3:0] _T_227; // @[LZD.scala 43:32]
  wire [1:0] _T_228; // @[LZD.scala 43:32]
  wire  _T_229; // @[LZD.scala 39:14]
  wire  _T_230; // @[LZD.scala 39:21]
  wire  _T_231; // @[LZD.scala 39:30]
  wire  _T_232; // @[LZD.scala 39:27]
  wire  _T_233; // @[LZD.scala 39:25]
  wire [1:0] _T_234; // @[Cat.scala 29:58]
  wire [1:0] _T_235; // @[LZD.scala 44:32]
  wire  _T_236; // @[LZD.scala 39:14]
  wire  _T_237; // @[LZD.scala 39:21]
  wire  _T_238; // @[LZD.scala 39:30]
  wire  _T_239; // @[LZD.scala 39:27]
  wire  _T_240; // @[LZD.scala 39:25]
  wire [1:0] _T_241; // @[Cat.scala 29:58]
  wire  _T_242; // @[Shift.scala 12:21]
  wire  _T_243; // @[Shift.scala 12:21]
  wire  _T_244; // @[LZD.scala 49:16]
  wire  _T_245; // @[LZD.scala 49:27]
  wire  _T_246; // @[LZD.scala 49:25]
  wire  _T_247; // @[LZD.scala 49:47]
  wire  _T_248; // @[LZD.scala 49:59]
  wire  _T_249; // @[LZD.scala 49:35]
  wire [2:0] _T_251; // @[Cat.scala 29:58]
  wire  _T_252; // @[LZD.scala 44:32]
  wire  _T_254; // @[Shift.scala 12:21]
  wire [1:0] _T_256; // @[Cat.scala 29:58]
  wire [1:0] _T_257; // @[LZD.scala 55:32]
  wire [1:0] _T_258; // @[LZD.scala 55:20]
  wire [2:0] _T_259; // @[Cat.scala 29:58]
  wire  _T_260; // @[Shift.scala 12:21]
  wire [2:0] _T_262; // @[LZD.scala 55:32]
  wire [2:0] _T_263; // @[LZD.scala 55:20]
  wire [3:0] _T_264; // @[Cat.scala 29:58]
  wire [3:0] _T_265; // @[convert.scala 21:22]
  wire [11:0] _T_266; // @[convert.scala 22:36]
  wire  _T_267; // @[Shift.scala 16:24]
  wire  _T_269; // @[Shift.scala 12:21]
  wire [3:0] _T_270; // @[Shift.scala 64:52]
  wire [11:0] _T_272; // @[Cat.scala 29:58]
  wire [11:0] _T_273; // @[Shift.scala 64:27]
  wire [2:0] _T_274; // @[Shift.scala 66:70]
  wire  _T_275; // @[Shift.scala 12:21]
  wire [7:0] _T_276; // @[Shift.scala 64:52]
  wire [11:0] _T_278; // @[Cat.scala 29:58]
  wire [11:0] _T_279; // @[Shift.scala 64:27]
  wire [1:0] _T_280; // @[Shift.scala 66:70]
  wire  _T_281; // @[Shift.scala 12:21]
  wire [9:0] _T_282; // @[Shift.scala 64:52]
  wire [11:0] _T_284; // @[Cat.scala 29:58]
  wire [11:0] _T_285; // @[Shift.scala 64:27]
  wire  _T_286; // @[Shift.scala 66:70]
  wire [10:0] _T_288; // @[Shift.scala 64:52]
  wire [11:0] _T_289; // @[Cat.scala 29:58]
  wire [11:0] _T_290; // @[Shift.scala 64:27]
  wire [11:0] _T_291; // @[Shift.scala 16:10]
  wire  _T_292; // @[convert.scala 23:34]
  wire [10:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_294; // @[convert.scala 25:26]
  wire [3:0] _T_296; // @[convert.scala 25:42]
  wire  _T_299; // @[convert.scala 26:67]
  wire  _T_300; // @[convert.scala 26:51]
  wire [5:0] _T_301; // @[Cat.scala 29:58]
  wire [13:0] _T_303; // @[convert.scala 29:56]
  wire  _T_304; // @[convert.scala 29:60]
  wire  _T_305; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_308; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_317; // @[Bitwise.scala 71:12]
  wire  _T_318; // @[PositDivisionSqrt.scala 80:40]
  wire [14:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_320; // @[PositDivisionSqrt.scala 82:31]
  wire [14:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_323; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_324; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_325; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_326; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_327; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_328; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_329; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_330; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_331; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_332; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [6:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_335; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_336; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_337; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_338; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_339; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_340; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_341; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_342; // @[PositDivisionSqrt.scala 117:30]
  wire [3:0] _T_344; // @[PositDivisionSqrt.scala 119:26]
  wire [3:0] _T_345; // @[PositDivisionSqrt.scala 118:20]
  wire [3:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [3:0] _T_346; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_348; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_349; // @[PositDivisionSqrt.scala 123:27]
  wire [3:0] _T_351; // @[PositDivisionSqrt.scala 123:52]
  wire [3:0] _T_352; // @[PositDivisionSqrt.scala 123:20]
  wire [3:0] _T_353; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_355; // @[PositDivisionSqrt.scala 124:27]
  wire [3:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_357; // @[PositDivisionSqrt.scala 123:64]
  wire [4:0] _T_358; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_360; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_361; // @[PositDivisionSqrt.scala 137:28]
  wire [15:0] _T_362; // @[PositDivisionSqrt.scala 146:22]
  wire [13:0] bitMask; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_364; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_365; // @[PositDivisionSqrt.scala 148:23]
  wire [14:0] _T_366; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_367; // @[PositDivisionSqrt.scala 149:23]
  wire [15:0] _T_368; // @[PositDivisionSqrt.scala 149:46]
  wire [14:0] _T_369; // @[PositDivisionSqrt.scala 149:56]
  wire [14:0] _T_370; // @[PositDivisionSqrt.scala 149:16]
  wire [14:0] _T_371; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_372; // @[PositDivisionSqrt.scala 150:17]
  wire [14:0] _T_373; // @[PositDivisionSqrt.scala 150:16]
  wire [14:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_375; // @[PositDivisionSqrt.scala 152:29]
  wire [14:0] _T_376; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_377; // @[PositDivisionSqrt.scala 153:29]
  wire [11:0] _T_378; // @[PositDivisionSqrt.scala 153:22]
  wire [14:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [14:0] _T_379; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_381; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_382; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_383; // @[PositDivisionSqrt.scala 154:57]
  wire [14:0] _T_386; // @[Cat.scala 29:58]
  wire [14:0] _T_387; // @[PositDivisionSqrt.scala 154:22]
  wire [14:0] _T_388; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_390; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_391; // @[PositDivisionSqrt.scala 156:79]
  wire [10:0] _T_393; // @[Bitwise.scala 71:12]
  wire [13:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [13:0] _T_394; // @[PositDivisionSqrt.scala 156:53]
  wire [14:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [14:0] _T_395; // @[PositDivisionSqrt.scala 155:51]
  wire [12:0] _T_396; // @[PositDivisionSqrt.scala 157:53]
  wire [14:0] _GEN_14; // @[PositDivisionSqrt.scala 156:85]
  wire [14:0] _T_397; // @[PositDivisionSqrt.scala 156:85]
  wire [14:0] _T_398; // @[PositDivisionSqrt.scala 155:22]
  wire [14:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_400; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_401; // @[PositDivisionSqrt.scala 162:40]
  wire [14:0] _T_404; // @[PositDivisionSqrt.scala 163:97]
  wire [14:0] _T_406; // @[PositDivisionSqrt.scala 164:97]
  wire [14:0] _T_407; // @[PositDivisionSqrt.scala 161:92]
  wire [15:0] _T_412; // @[PositDivisionSqrt.scala 168:98]
  wire [14:0] _T_413; // @[PositDivisionSqrt.scala 168:108]
  wire [14:0] _T_415; // @[PositDivisionSqrt.scala 168:112]
  wire [14:0] _T_419; // @[PositDivisionSqrt.scala 169:112]
  wire [14:0] _T_420; // @[PositDivisionSqrt.scala 166:26]
  wire [14:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_421; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_422; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_424; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_425; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_426; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_427; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_428; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_430; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_431; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_432; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_433; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_434; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_437; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_438; // @[PositDivisionSqrt.scala 187:28]
  wire [14:0] _T_441; // @[PositDivisionSqrt.scala 188:47]
  wire [14:0] _T_442; // @[PositDivisionSqrt.scala 188:18]
  wire [12:0] _T_444; // @[PositDivisionSqrt.scala 189:18]
  wire [14:0] _GEN_15; // @[PositDivisionSqrt.scala 188:72]
  wire [14:0] _T_445; // @[PositDivisionSqrt.scala 188:72]
  wire [14:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [14:0] _T_447; // @[PositDivisionSqrt.scala 190:47]
  wire [14:0] _T_448; // @[PositDivisionSqrt.scala 190:18]
  wire [14:0] _T_449; // @[PositDivisionSqrt.scala 189:72]
  wire [1:0] _T_451; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [14:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [14:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [10:0] _T_454; // @[PositDivisionSqrt.scala 200:97]
  wire [10:0] _T_455; // @[PositDivisionSqrt.scala 201:97]
  wire [10:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_456; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_457; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_458; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_460; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_461; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_462; // @[Cat.scala 29:58]
  wire [2:0] _T_463; // @[PositDivisionSqrt.scala 209:63]
  wire [6:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] _T_465; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [6:0] _T_467; // @[Mux.scala 87:16]
  wire [6:0] _T_468; // @[Mux.scala 87:16]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [5:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [5:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire  _T_473; // @[convert.scala 46:61]
  wire  _T_474; // @[convert.scala 46:52]
  wire  _T_476; // @[convert.scala 46:42]
  wire [4:0] _T_477; // @[convert.scala 48:34]
  wire  _T_478; // @[convert.scala 49:36]
  wire [4:0] _T_480; // @[convert.scala 50:36]
  wire [4:0] _T_481; // @[convert.scala 50:36]
  wire [4:0] _T_482; // @[convert.scala 50:28]
  wire  _T_483; // @[convert.scala 51:31]
  wire  _T_484; // @[convert.scala 52:43]
  wire [16:0] _T_488; // @[Cat.scala 29:58]
  wire [4:0] _T_489; // @[Shift.scala 39:17]
  wire  _T_490; // @[Shift.scala 39:24]
  wire  _T_492; // @[Shift.scala 90:30]
  wire [15:0] _T_493; // @[Shift.scala 90:48]
  wire  _T_494; // @[Shift.scala 90:57]
  wire  _T_495; // @[Shift.scala 90:39]
  wire  _T_496; // @[Shift.scala 12:21]
  wire  _T_497; // @[Shift.scala 12:21]
  wire [15:0] _T_499; // @[Bitwise.scala 71:12]
  wire [16:0] _T_500; // @[Cat.scala 29:58]
  wire [16:0] _T_501; // @[Shift.scala 91:22]
  wire [3:0] _T_502; // @[Shift.scala 92:77]
  wire [8:0] _T_503; // @[Shift.scala 90:30]
  wire [7:0] _T_504; // @[Shift.scala 90:48]
  wire  _T_505; // @[Shift.scala 90:57]
  wire [8:0] _GEN_20; // @[Shift.scala 90:39]
  wire [8:0] _T_506; // @[Shift.scala 90:39]
  wire  _T_507; // @[Shift.scala 12:21]
  wire  _T_508; // @[Shift.scala 12:21]
  wire [7:0] _T_510; // @[Bitwise.scala 71:12]
  wire [16:0] _T_511; // @[Cat.scala 29:58]
  wire [16:0] _T_512; // @[Shift.scala 91:22]
  wire [2:0] _T_513; // @[Shift.scala 92:77]
  wire [12:0] _T_514; // @[Shift.scala 90:30]
  wire [3:0] _T_515; // @[Shift.scala 90:48]
  wire  _T_516; // @[Shift.scala 90:57]
  wire [12:0] _GEN_21; // @[Shift.scala 90:39]
  wire [12:0] _T_517; // @[Shift.scala 90:39]
  wire  _T_518; // @[Shift.scala 12:21]
  wire  _T_519; // @[Shift.scala 12:21]
  wire [3:0] _T_521; // @[Bitwise.scala 71:12]
  wire [16:0] _T_522; // @[Cat.scala 29:58]
  wire [16:0] _T_523; // @[Shift.scala 91:22]
  wire [1:0] _T_524; // @[Shift.scala 92:77]
  wire [14:0] _T_525; // @[Shift.scala 90:30]
  wire [1:0] _T_526; // @[Shift.scala 90:48]
  wire  _T_527; // @[Shift.scala 90:57]
  wire [14:0] _GEN_22; // @[Shift.scala 90:39]
  wire [14:0] _T_528; // @[Shift.scala 90:39]
  wire  _T_529; // @[Shift.scala 12:21]
  wire  _T_530; // @[Shift.scala 12:21]
  wire [1:0] _T_532; // @[Bitwise.scala 71:12]
  wire [16:0] _T_533; // @[Cat.scala 29:58]
  wire [16:0] _T_534; // @[Shift.scala 91:22]
  wire  _T_535; // @[Shift.scala 92:77]
  wire [15:0] _T_536; // @[Shift.scala 90:30]
  wire  _T_537; // @[Shift.scala 90:48]
  wire [15:0] _GEN_23; // @[Shift.scala 90:39]
  wire [15:0] _T_539; // @[Shift.scala 90:39]
  wire  _T_541; // @[Shift.scala 12:21]
  wire [16:0] _T_542; // @[Cat.scala 29:58]
  wire [16:0] _T_543; // @[Shift.scala 91:22]
  wire [16:0] _T_546; // @[Bitwise.scala 71:12]
  wire [16:0] _T_547; // @[Shift.scala 39:10]
  wire  _T_548; // @[convert.scala 55:31]
  wire  _T_549; // @[convert.scala 56:31]
  wire  _T_550; // @[convert.scala 57:31]
  wire  _T_551; // @[convert.scala 58:31]
  wire [13:0] _T_552; // @[convert.scala 59:69]
  wire  _T_553; // @[convert.scala 59:81]
  wire  _T_554; // @[convert.scala 59:50]
  wire  _T_556; // @[convert.scala 60:81]
  wire  _T_557; // @[convert.scala 61:44]
  wire  _T_558; // @[convert.scala 61:52]
  wire  _T_559; // @[convert.scala 61:36]
  wire  _T_560; // @[convert.scala 62:63]
  wire  _T_561; // @[convert.scala 62:103]
  wire  _T_562; // @[convert.scala 62:60]
  wire [13:0] _GEN_24; // @[convert.scala 63:56]
  wire [13:0] _T_565; // @[convert.scala 63:56]
  wire [14:0] _T_566; // @[Cat.scala 29:58]
  wire [14:0] _T_568; // @[Mux.scala 87:16]
  assign _T_1 = io_A[14]; // @[convert.scala 18:24]
  assign _T_2 = io_A[13]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[13:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[12:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[12:5]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[4:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68[4:1]; // @[LZD.scala 43:32]
  assign _T_70 = _T_69[3:2]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70 != 2'h0; // @[LZD.scala 39:14]
  assign _T_72 = _T_70[1]; // @[LZD.scala 39:21]
  assign _T_73 = _T_70[0]; // @[LZD.scala 39:30]
  assign _T_74 = ~ _T_73; // @[LZD.scala 39:27]
  assign _T_75 = _T_72 | _T_74; // @[LZD.scala 39:25]
  assign _T_76 = {_T_71,_T_75}; // @[Cat.scala 29:58]
  assign _T_77 = _T_69[1:0]; // @[LZD.scala 44:32]
  assign _T_78 = _T_77 != 2'h0; // @[LZD.scala 39:14]
  assign _T_79 = _T_77[1]; // @[LZD.scala 39:21]
  assign _T_80 = _T_77[0]; // @[LZD.scala 39:30]
  assign _T_81 = ~ _T_80; // @[LZD.scala 39:27]
  assign _T_82 = _T_79 | _T_81; // @[LZD.scala 39:25]
  assign _T_83 = {_T_78,_T_82}; // @[Cat.scala 29:58]
  assign _T_84 = _T_76[1]; // @[Shift.scala 12:21]
  assign _T_85 = _T_83[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84 | _T_85; // @[LZD.scala 49:16]
  assign _T_87 = ~ _T_85; // @[LZD.scala 49:27]
  assign _T_88 = _T_84 | _T_87; // @[LZD.scala 49:25]
  assign _T_89 = _T_76[0:0]; // @[LZD.scala 49:47]
  assign _T_90 = _T_83[0:0]; // @[LZD.scala 49:59]
  assign _T_91 = _T_84 ? _T_89 : _T_90; // @[LZD.scala 49:35]
  assign _T_93 = {_T_86,_T_88,_T_91}; // @[Cat.scala 29:58]
  assign _T_94 = _T_68[0:0]; // @[LZD.scala 44:32]
  assign _T_96 = _T_93[2]; // @[Shift.scala 12:21]
  assign _T_98 = {1'h1,_T_94}; // @[Cat.scala 29:58]
  assign _T_99 = _T_93[1:0]; // @[LZD.scala 55:32]
  assign _T_100 = _T_96 ? _T_99 : _T_98; // @[LZD.scala 55:20]
  assign _T_101 = {_T_96,_T_100}; // @[Cat.scala 29:58]
  assign _T_102 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_104 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_105 = _T_102 ? _T_104 : _T_101; // @[LZD.scala 55:20]
  assign _T_106 = {_T_102,_T_105}; // @[Cat.scala 29:58]
  assign _T_107 = ~ _T_106; // @[convert.scala 21:22]
  assign _T_108 = io_A[11:0]; // @[convert.scala 22:36]
  assign _T_109 = _T_107 < 4'hc; // @[Shift.scala 16:24]
  assign _T_111 = _T_107[3]; // @[Shift.scala 12:21]
  assign _T_112 = _T_108[3:0]; // @[Shift.scala 64:52]
  assign _T_114 = {_T_112,8'h0}; // @[Cat.scala 29:58]
  assign _T_115 = _T_111 ? _T_114 : _T_108; // @[Shift.scala 64:27]
  assign _T_116 = _T_107[2:0]; // @[Shift.scala 66:70]
  assign _T_117 = _T_116[2]; // @[Shift.scala 12:21]
  assign _T_118 = _T_115[7:0]; // @[Shift.scala 64:52]
  assign _T_120 = {_T_118,4'h0}; // @[Cat.scala 29:58]
  assign _T_121 = _T_117 ? _T_120 : _T_115; // @[Shift.scala 64:27]
  assign _T_122 = _T_116[1:0]; // @[Shift.scala 66:70]
  assign _T_123 = _T_122[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_121[9:0]; // @[Shift.scala 64:52]
  assign _T_126 = {_T_124,2'h0}; // @[Cat.scala 29:58]
  assign _T_127 = _T_123 ? _T_126 : _T_121; // @[Shift.scala 64:27]
  assign _T_128 = _T_122[0:0]; // @[Shift.scala 66:70]
  assign _T_130 = _T_127[10:0]; // @[Shift.scala 64:52]
  assign _T_131 = {_T_130,1'h0}; // @[Cat.scala 29:58]
  assign _T_132 = _T_128 ? _T_131 : _T_127; // @[Shift.scala 64:27]
  assign _T_133 = _T_109 ? _T_132 : 12'h0; // @[Shift.scala 16:10]
  assign _T_134 = _T_133[11:11]; // @[convert.scala 23:34]
  assign decA_fraction = _T_133[10:0]; // @[convert.scala 24:34]
  assign _T_136 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_138 = _T_3 ? _T_107 : _T_106; // @[convert.scala 25:42]
  assign _T_141 = ~ _T_134; // @[convert.scala 26:67]
  assign _T_142 = _T_1 ? _T_141 : _T_134; // @[convert.scala 26:51]
  assign _T_143 = {_T_136,_T_138,_T_142}; // @[Cat.scala 29:58]
  assign _T_145 = io_A[13:0]; // @[convert.scala 29:56]
  assign _T_146 = _T_145 != 14'h0; // @[convert.scala 29:60]
  assign _T_147 = ~ _T_146; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_147; // @[convert.scala 29:39]
  assign _T_150 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_150 & _T_147; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_143); // @[convert.scala 32:24]
  assign _T_159 = io_B[14]; // @[convert.scala 18:24]
  assign _T_160 = io_B[13]; // @[convert.scala 18:40]
  assign _T_161 = _T_159 ^ _T_160; // @[convert.scala 18:36]
  assign _T_162 = io_B[13:1]; // @[convert.scala 19:24]
  assign _T_163 = io_B[12:0]; // @[convert.scala 19:43]
  assign _T_164 = _T_162 ^ _T_163; // @[convert.scala 19:39]
  assign _T_165 = _T_164[12:5]; // @[LZD.scala 43:32]
  assign _T_166 = _T_165[7:4]; // @[LZD.scala 43:32]
  assign _T_167 = _T_166[3:2]; // @[LZD.scala 43:32]
  assign _T_168 = _T_167 != 2'h0; // @[LZD.scala 39:14]
  assign _T_169 = _T_167[1]; // @[LZD.scala 39:21]
  assign _T_170 = _T_167[0]; // @[LZD.scala 39:30]
  assign _T_171 = ~ _T_170; // @[LZD.scala 39:27]
  assign _T_172 = _T_169 | _T_171; // @[LZD.scala 39:25]
  assign _T_173 = {_T_168,_T_172}; // @[Cat.scala 29:58]
  assign _T_174 = _T_166[1:0]; // @[LZD.scala 44:32]
  assign _T_175 = _T_174 != 2'h0; // @[LZD.scala 39:14]
  assign _T_176 = _T_174[1]; // @[LZD.scala 39:21]
  assign _T_177 = _T_174[0]; // @[LZD.scala 39:30]
  assign _T_178 = ~ _T_177; // @[LZD.scala 39:27]
  assign _T_179 = _T_176 | _T_178; // @[LZD.scala 39:25]
  assign _T_180 = {_T_175,_T_179}; // @[Cat.scala 29:58]
  assign _T_181 = _T_173[1]; // @[Shift.scala 12:21]
  assign _T_182 = _T_180[1]; // @[Shift.scala 12:21]
  assign _T_183 = _T_181 | _T_182; // @[LZD.scala 49:16]
  assign _T_184 = ~ _T_182; // @[LZD.scala 49:27]
  assign _T_185 = _T_181 | _T_184; // @[LZD.scala 49:25]
  assign _T_186 = _T_173[0:0]; // @[LZD.scala 49:47]
  assign _T_187 = _T_180[0:0]; // @[LZD.scala 49:59]
  assign _T_188 = _T_181 ? _T_186 : _T_187; // @[LZD.scala 49:35]
  assign _T_190 = {_T_183,_T_185,_T_188}; // @[Cat.scala 29:58]
  assign _T_191 = _T_165[3:0]; // @[LZD.scala 44:32]
  assign _T_192 = _T_191[3:2]; // @[LZD.scala 43:32]
  assign _T_193 = _T_192 != 2'h0; // @[LZD.scala 39:14]
  assign _T_194 = _T_192[1]; // @[LZD.scala 39:21]
  assign _T_195 = _T_192[0]; // @[LZD.scala 39:30]
  assign _T_196 = ~ _T_195; // @[LZD.scala 39:27]
  assign _T_197 = _T_194 | _T_196; // @[LZD.scala 39:25]
  assign _T_198 = {_T_193,_T_197}; // @[Cat.scala 29:58]
  assign _T_199 = _T_191[1:0]; // @[LZD.scala 44:32]
  assign _T_200 = _T_199 != 2'h0; // @[LZD.scala 39:14]
  assign _T_201 = _T_199[1]; // @[LZD.scala 39:21]
  assign _T_202 = _T_199[0]; // @[LZD.scala 39:30]
  assign _T_203 = ~ _T_202; // @[LZD.scala 39:27]
  assign _T_204 = _T_201 | _T_203; // @[LZD.scala 39:25]
  assign _T_205 = {_T_200,_T_204}; // @[Cat.scala 29:58]
  assign _T_206 = _T_198[1]; // @[Shift.scala 12:21]
  assign _T_207 = _T_205[1]; // @[Shift.scala 12:21]
  assign _T_208 = _T_206 | _T_207; // @[LZD.scala 49:16]
  assign _T_209 = ~ _T_207; // @[LZD.scala 49:27]
  assign _T_210 = _T_206 | _T_209; // @[LZD.scala 49:25]
  assign _T_211 = _T_198[0:0]; // @[LZD.scala 49:47]
  assign _T_212 = _T_205[0:0]; // @[LZD.scala 49:59]
  assign _T_213 = _T_206 ? _T_211 : _T_212; // @[LZD.scala 49:35]
  assign _T_215 = {_T_208,_T_210,_T_213}; // @[Cat.scala 29:58]
  assign _T_216 = _T_190[2]; // @[Shift.scala 12:21]
  assign _T_217 = _T_215[2]; // @[Shift.scala 12:21]
  assign _T_218 = _T_216 | _T_217; // @[LZD.scala 49:16]
  assign _T_219 = ~ _T_217; // @[LZD.scala 49:27]
  assign _T_220 = _T_216 | _T_219; // @[LZD.scala 49:25]
  assign _T_221 = _T_190[1:0]; // @[LZD.scala 49:47]
  assign _T_222 = _T_215[1:0]; // @[LZD.scala 49:59]
  assign _T_223 = _T_216 ? _T_221 : _T_222; // @[LZD.scala 49:35]
  assign _T_225 = {_T_218,_T_220,_T_223}; // @[Cat.scala 29:58]
  assign _T_226 = _T_164[4:0]; // @[LZD.scala 44:32]
  assign _T_227 = _T_226[4:1]; // @[LZD.scala 43:32]
  assign _T_228 = _T_227[3:2]; // @[LZD.scala 43:32]
  assign _T_229 = _T_228 != 2'h0; // @[LZD.scala 39:14]
  assign _T_230 = _T_228[1]; // @[LZD.scala 39:21]
  assign _T_231 = _T_228[0]; // @[LZD.scala 39:30]
  assign _T_232 = ~ _T_231; // @[LZD.scala 39:27]
  assign _T_233 = _T_230 | _T_232; // @[LZD.scala 39:25]
  assign _T_234 = {_T_229,_T_233}; // @[Cat.scala 29:58]
  assign _T_235 = _T_227[1:0]; // @[LZD.scala 44:32]
  assign _T_236 = _T_235 != 2'h0; // @[LZD.scala 39:14]
  assign _T_237 = _T_235[1]; // @[LZD.scala 39:21]
  assign _T_238 = _T_235[0]; // @[LZD.scala 39:30]
  assign _T_239 = ~ _T_238; // @[LZD.scala 39:27]
  assign _T_240 = _T_237 | _T_239; // @[LZD.scala 39:25]
  assign _T_241 = {_T_236,_T_240}; // @[Cat.scala 29:58]
  assign _T_242 = _T_234[1]; // @[Shift.scala 12:21]
  assign _T_243 = _T_241[1]; // @[Shift.scala 12:21]
  assign _T_244 = _T_242 | _T_243; // @[LZD.scala 49:16]
  assign _T_245 = ~ _T_243; // @[LZD.scala 49:27]
  assign _T_246 = _T_242 | _T_245; // @[LZD.scala 49:25]
  assign _T_247 = _T_234[0:0]; // @[LZD.scala 49:47]
  assign _T_248 = _T_241[0:0]; // @[LZD.scala 49:59]
  assign _T_249 = _T_242 ? _T_247 : _T_248; // @[LZD.scala 49:35]
  assign _T_251 = {_T_244,_T_246,_T_249}; // @[Cat.scala 29:58]
  assign _T_252 = _T_226[0:0]; // @[LZD.scala 44:32]
  assign _T_254 = _T_251[2]; // @[Shift.scala 12:21]
  assign _T_256 = {1'h1,_T_252}; // @[Cat.scala 29:58]
  assign _T_257 = _T_251[1:0]; // @[LZD.scala 55:32]
  assign _T_258 = _T_254 ? _T_257 : _T_256; // @[LZD.scala 55:20]
  assign _T_259 = {_T_254,_T_258}; // @[Cat.scala 29:58]
  assign _T_260 = _T_225[3]; // @[Shift.scala 12:21]
  assign _T_262 = _T_225[2:0]; // @[LZD.scala 55:32]
  assign _T_263 = _T_260 ? _T_262 : _T_259; // @[LZD.scala 55:20]
  assign _T_264 = {_T_260,_T_263}; // @[Cat.scala 29:58]
  assign _T_265 = ~ _T_264; // @[convert.scala 21:22]
  assign _T_266 = io_B[11:0]; // @[convert.scala 22:36]
  assign _T_267 = _T_265 < 4'hc; // @[Shift.scala 16:24]
  assign _T_269 = _T_265[3]; // @[Shift.scala 12:21]
  assign _T_270 = _T_266[3:0]; // @[Shift.scala 64:52]
  assign _T_272 = {_T_270,8'h0}; // @[Cat.scala 29:58]
  assign _T_273 = _T_269 ? _T_272 : _T_266; // @[Shift.scala 64:27]
  assign _T_274 = _T_265[2:0]; // @[Shift.scala 66:70]
  assign _T_275 = _T_274[2]; // @[Shift.scala 12:21]
  assign _T_276 = _T_273[7:0]; // @[Shift.scala 64:52]
  assign _T_278 = {_T_276,4'h0}; // @[Cat.scala 29:58]
  assign _T_279 = _T_275 ? _T_278 : _T_273; // @[Shift.scala 64:27]
  assign _T_280 = _T_274[1:0]; // @[Shift.scala 66:70]
  assign _T_281 = _T_280[1]; // @[Shift.scala 12:21]
  assign _T_282 = _T_279[9:0]; // @[Shift.scala 64:52]
  assign _T_284 = {_T_282,2'h0}; // @[Cat.scala 29:58]
  assign _T_285 = _T_281 ? _T_284 : _T_279; // @[Shift.scala 64:27]
  assign _T_286 = _T_280[0:0]; // @[Shift.scala 66:70]
  assign _T_288 = _T_285[10:0]; // @[Shift.scala 64:52]
  assign _T_289 = {_T_288,1'h0}; // @[Cat.scala 29:58]
  assign _T_290 = _T_286 ? _T_289 : _T_285; // @[Shift.scala 64:27]
  assign _T_291 = _T_267 ? _T_290 : 12'h0; // @[Shift.scala 16:10]
  assign _T_292 = _T_291[11:11]; // @[convert.scala 23:34]
  assign decB_fraction = _T_291[10:0]; // @[convert.scala 24:34]
  assign _T_294 = _T_161 == 1'h0; // @[convert.scala 25:26]
  assign _T_296 = _T_161 ? _T_265 : _T_264; // @[convert.scala 25:42]
  assign _T_299 = ~ _T_292; // @[convert.scala 26:67]
  assign _T_300 = _T_159 ? _T_299 : _T_292; // @[convert.scala 26:51]
  assign _T_301 = {_T_294,_T_296,_T_300}; // @[Cat.scala 29:58]
  assign _T_303 = io_B[13:0]; // @[convert.scala 29:56]
  assign _T_304 = _T_303 != 14'h0; // @[convert.scala 29:60]
  assign _T_305 = ~ _T_304; // @[convert.scala 29:41]
  assign decB_isNaR = _T_159 & _T_305; // @[convert.scala 29:39]
  assign _T_308 = _T_159 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_308 & _T_305; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_301); // @[convert.scala 32:24]
  assign _T_317 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_318 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_317,_T_318,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_320 = ~ _T_159; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_159,_T_320,decB_fraction,2'h0}; // @[Cat.scala 29:58]
  assign _T_323 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_323 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_324 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_325 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_326 = _T_325 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_327 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_328 = decA_isZero & _T_327; // @[PositDivisionSqrt.scala 94:43]
  assign _T_329 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_330 = _T_328 & _T_329; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_331 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_332 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_331 & _T_332; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_331 & _T_150; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_335 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_335; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 4'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_336 = sigX_Z[14]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_337 = sigX_Z[12]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_336 ^ _T_337; // @[PositDivisionSqrt.scala 113:50]
  assign _T_338 = cycleNum == 4'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_338 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_339 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_340 = _T_339 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_341 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_342 = entering & _T_341; // @[PositDivisionSqrt.scala 117:30]
  assign _T_344 = io_sqrtOp ? 4'hd : 4'hf; // @[PositDivisionSqrt.scala 119:26]
  assign _T_345 = entering_normalCase ? _T_344 : 4'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{3'd0}, _T_342}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_346 = _GEN_9 | _T_345; // @[PositDivisionSqrt.scala 117:64]
  assign _T_348 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_349 = _T_339 & _T_348; // @[PositDivisionSqrt.scala 123:27]
  assign _T_351 = cycleNum - 4'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_352 = _T_349 ? _T_351 : 4'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_353 = _T_346 | _T_352; // @[PositDivisionSqrt.scala 122:64]
  assign _T_355 = _T_339 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{3'd0}, _T_355}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_357 = _T_353 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_358 = decA_scale[5:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_360 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_361 = entering_normalCase & _T_360; // @[PositDivisionSqrt.scala 137:28]
  assign _T_362 = 16'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign bitMask = _T_362[15:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_364 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_365 = ready & _T_364; // @[PositDivisionSqrt.scala 148:23]
  assign _T_366 = _T_365 ? sigA_S : 15'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_367 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_368 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_369 = _T_368[14:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_370 = _T_367 ? _T_369 : 15'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_371 = _T_366 | _T_370; // @[PositDivisionSqrt.scala 148:66]
  assign _T_372 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_373 = _T_372 ? rem_Z : 15'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_371 | _T_373; // @[PositDivisionSqrt.scala 149:66]
  assign _T_375 = ready & _T_360; // @[PositDivisionSqrt.scala 152:29]
  assign _T_376 = _T_375 ? sigB_S : 15'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_377 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_378 = _T_377 ? 12'h800 : 12'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_378}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_379 = _T_376 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_381 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_382 = _T_372 & _T_381; // @[PositDivisionSqrt.scala 154:30]
  assign _T_383 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_386 = {signB_Z,_T_383,fractB_Z,2'h0}; // @[Cat.scala 29:58]
  assign _T_387 = _T_382 ? _T_386 : 15'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_388 = _T_379 | _T_387; // @[PositDivisionSqrt.scala 153:93]
  assign _T_390 = _T_372 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_391 = rem[14:14]; // @[PositDivisionSqrt.scala 156:79]
  assign _T_393 = _T_391 ? 11'h7ff : 11'h0; // @[Bitwise.scala 71:12]
  assign _GEN_12 = {{3'd0}, _T_393}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_394 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_394}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_395 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_396 = bitMask[13:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_396}; // @[PositDivisionSqrt.scala 156:85]
  assign _T_397 = _T_395 | _GEN_14; // @[PositDivisionSqrt.scala 156:85]
  assign _T_398 = _T_390 ? _T_397 : 15'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_388 | _T_398; // @[PositDivisionSqrt.scala 154:93]
  assign _T_400 = trialTerm[14:14]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_401 = _T_391 ^ _T_400; // @[PositDivisionSqrt.scala 162:40]
  assign _T_404 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_406 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_407 = _T_401 ? _T_404 : _T_406; // @[PositDivisionSqrt.scala 161:92]
  assign _T_412 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_413 = _T_412[14:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_415 = _T_413 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_419 = _T_413 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_420 = _T_401 ? _T_415 : _T_419; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_407 : _T_420; // @[PositDivisionSqrt.scala 159:27]
  assign _T_421 = trialRem != 15'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_421 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_422 = rem != 15'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_422 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_424 = trialRem[14:14]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_425 = _T_400 ^ _T_424; // @[PositDivisionSqrt.scala 176:49]
  assign _T_426 = ~ _T_425; // @[PositDivisionSqrt.scala 176:29]
  assign _T_427 = sigX_Z[14:14]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_428 = ~ _T_427; // @[PositDivisionSqrt.scala 178:49]
  assign _T_430 = remIsZero ? _T_427 : _T_426; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_428 : _T_430; // @[Mux.scala 87:16]
  assign _T_431 = cycleNum > 4'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_432 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_433 = _T_431 & _T_432; // @[PositDivisionSqrt.scala 183:48]
  assign _T_434 = entering_normalCase | _T_433; // @[PositDivisionSqrt.scala 183:28]
  assign _T_437 = _T_372 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_438 = entering_normalCase | _T_437; // @[PositDivisionSqrt.scala 187:28]
  assign _T_441 = {newBit, 14'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_442 = _T_375 ? _T_441 : 15'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_444 = _T_377 ? 13'h1000 : 13'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_444}; // @[PositDivisionSqrt.scala 188:72]
  assign _T_445 = _T_442 | _GEN_15; // @[PositDivisionSqrt.scala 188:72]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_447 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_448 = _T_372 ? _T_447 : 15'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_449 = _T_445 | _T_448; // @[PositDivisionSqrt.scala 189:72]
  assign _T_451 = {_T_427, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_451 : {{1'd0}, _T_427}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{13'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_454 = realSigX[11:1]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_455 = realSigX[10:0]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_454 : _T_455; // @[PositDivisionSqrt.scala 198:21]
  assign _T_456 = realSigX[14]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_457 = realSigX[12]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_458 = _T_456 ^ _T_457; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_458; // @[PositDivisionSqrt.scala 205:23]
  assign _T_460 = realSigX[11]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_456 ^ _T_460; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_461 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_461; // @[PositDivisionSqrt.scala 208:36]
  assign _T_462 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_463 = {1'b0,$signed(_T_462)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{4{_T_463[2]}},_T_463}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_465 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_465); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-7'sh1a); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(7'sh1a); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[14:14]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_467 = underflow ? $signed(-7'sh1a) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_468 = overflow ? $signed(7'sh1a) : $signed(_T_467); // @[Mux.scala 87:16]
  assign outValid = cycleNum == 4'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_468[5:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_473 = decQ_scale[0]; // @[convert.scala 46:61]
  assign _T_474 = ~ _T_473; // @[convert.scala 46:52]
  assign _T_476 = decQ_sign ? _T_474 : _T_473; // @[convert.scala 46:42]
  assign _T_477 = decQ_scale[5:1]; // @[convert.scala 48:34]
  assign _T_478 = _T_477[4:4]; // @[convert.scala 49:36]
  assign _T_480 = ~ _T_477; // @[convert.scala 50:36]
  assign _T_481 = $signed(_T_480); // @[convert.scala 50:36]
  assign _T_482 = _T_478 ? $signed(_T_481) : $signed(_T_477); // @[convert.scala 50:28]
  assign _T_483 = _T_478 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_484 = ~ _T_483; // @[convert.scala 52:43]
  assign _T_488 = {_T_484,_T_483,_T_476,realFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_489 = $unsigned(_T_482); // @[Shift.scala 39:17]
  assign _T_490 = _T_489 < 5'h11; // @[Shift.scala 39:24]
  assign _T_492 = _T_488[16:16]; // @[Shift.scala 90:30]
  assign _T_493 = _T_488[15:0]; // @[Shift.scala 90:48]
  assign _T_494 = _T_493 != 16'h0; // @[Shift.scala 90:57]
  assign _T_495 = _T_492 | _T_494; // @[Shift.scala 90:39]
  assign _T_496 = _T_489[4]; // @[Shift.scala 12:21]
  assign _T_497 = _T_488[16]; // @[Shift.scala 12:21]
  assign _T_499 = _T_497 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_500 = {_T_499,_T_495}; // @[Cat.scala 29:58]
  assign _T_501 = _T_496 ? _T_500 : _T_488; // @[Shift.scala 91:22]
  assign _T_502 = _T_489[3:0]; // @[Shift.scala 92:77]
  assign _T_503 = _T_501[16:8]; // @[Shift.scala 90:30]
  assign _T_504 = _T_501[7:0]; // @[Shift.scala 90:48]
  assign _T_505 = _T_504 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{8'd0}, _T_505}; // @[Shift.scala 90:39]
  assign _T_506 = _T_503 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_507 = _T_502[3]; // @[Shift.scala 12:21]
  assign _T_508 = _T_501[16]; // @[Shift.scala 12:21]
  assign _T_510 = _T_508 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_511 = {_T_510,_T_506}; // @[Cat.scala 29:58]
  assign _T_512 = _T_507 ? _T_511 : _T_501; // @[Shift.scala 91:22]
  assign _T_513 = _T_502[2:0]; // @[Shift.scala 92:77]
  assign _T_514 = _T_512[16:4]; // @[Shift.scala 90:30]
  assign _T_515 = _T_512[3:0]; // @[Shift.scala 90:48]
  assign _T_516 = _T_515 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{12'd0}, _T_516}; // @[Shift.scala 90:39]
  assign _T_517 = _T_514 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_518 = _T_513[2]; // @[Shift.scala 12:21]
  assign _T_519 = _T_512[16]; // @[Shift.scala 12:21]
  assign _T_521 = _T_519 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_522 = {_T_521,_T_517}; // @[Cat.scala 29:58]
  assign _T_523 = _T_518 ? _T_522 : _T_512; // @[Shift.scala 91:22]
  assign _T_524 = _T_513[1:0]; // @[Shift.scala 92:77]
  assign _T_525 = _T_523[16:2]; // @[Shift.scala 90:30]
  assign _T_526 = _T_523[1:0]; // @[Shift.scala 90:48]
  assign _T_527 = _T_526 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{14'd0}, _T_527}; // @[Shift.scala 90:39]
  assign _T_528 = _T_525 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_529 = _T_524[1]; // @[Shift.scala 12:21]
  assign _T_530 = _T_523[16]; // @[Shift.scala 12:21]
  assign _T_532 = _T_530 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_533 = {_T_532,_T_528}; // @[Cat.scala 29:58]
  assign _T_534 = _T_529 ? _T_533 : _T_523; // @[Shift.scala 91:22]
  assign _T_535 = _T_524[0:0]; // @[Shift.scala 92:77]
  assign _T_536 = _T_534[16:1]; // @[Shift.scala 90:30]
  assign _T_537 = _T_534[0:0]; // @[Shift.scala 90:48]
  assign _GEN_23 = {{15'd0}, _T_537}; // @[Shift.scala 90:39]
  assign _T_539 = _T_536 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_541 = _T_534[16]; // @[Shift.scala 12:21]
  assign _T_542 = {_T_541,_T_539}; // @[Cat.scala 29:58]
  assign _T_543 = _T_535 ? _T_542 : _T_534; // @[Shift.scala 91:22]
  assign _T_546 = _T_497 ? 17'h1ffff : 17'h0; // @[Bitwise.scala 71:12]
  assign _T_547 = _T_490 ? _T_543 : _T_546; // @[Shift.scala 39:10]
  assign _T_548 = _T_547[3]; // @[convert.scala 55:31]
  assign _T_549 = _T_547[2]; // @[convert.scala 56:31]
  assign _T_550 = _T_547[1]; // @[convert.scala 57:31]
  assign _T_551 = _T_547[0]; // @[convert.scala 58:31]
  assign _T_552 = _T_547[16:3]; // @[convert.scala 59:69]
  assign _T_553 = _T_552 != 14'h0; // @[convert.scala 59:81]
  assign _T_554 = ~ _T_553; // @[convert.scala 59:50]
  assign _T_556 = _T_552 == 14'h3fff; // @[convert.scala 60:81]
  assign _T_557 = _T_548 | _T_550; // @[convert.scala 61:44]
  assign _T_558 = _T_557 | _T_551; // @[convert.scala 61:52]
  assign _T_559 = _T_549 & _T_558; // @[convert.scala 61:36]
  assign _T_560 = ~ _T_556; // @[convert.scala 62:63]
  assign _T_561 = _T_560 & _T_559; // @[convert.scala 62:103]
  assign _T_562 = _T_554 | _T_561; // @[convert.scala 62:60]
  assign _GEN_24 = {{13'd0}, _T_562}; // @[convert.scala 63:56]
  assign _T_565 = _T_552 + _GEN_24; // @[convert.scala 63:56]
  assign _T_566 = {decQ_sign,_T_565}; // @[Cat.scala 29:58]
  assign _T_568 = isZero_Z ? 15'h0 : _T_566; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_381; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 15'h4000 : _T_568; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[14:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 4'h0;
    end else begin
      if (_T_340) begin
        cycleNum <= _T_357;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_324;
      end else begin
        isNaR_Z <= _T_326;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_330;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_358[4]}},_T_358};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_361) begin
      signB_Z <= _T_159;
    end
    if (_T_361) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_434) begin
      if (ready) begin
        if (_T_401) begin
          rem_Z <= _T_404;
        end else begin
          rem_Z <= _T_406;
        end
      end else begin
        if (_T_401) begin
          rem_Z <= _T_415;
        end else begin
          rem_Z <= _T_419;
        end
      end
    end
    if (_T_438) begin
      sigX_Z <= _T_449;
    end
  end
endmodule
