module PositAdder29_3(
  input         clock,
  input         reset,
  input  [28:0] io_A,
  input  [28:0] io_B,
  output [28:0] io_S
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [26:0] _T_4; // @[convert.scala 19:24]
  wire [26:0] _T_5; // @[convert.scala 19:43]
  wire [26:0] _T_6; // @[convert.scala 19:39]
  wire [15:0] _T_7; // @[LZD.scala 43:32]
  wire [7:0] _T_8; // @[LZD.scala 43:32]
  wire [3:0] _T_9; // @[LZD.scala 43:32]
  wire [1:0] _T_10; // @[LZD.scala 43:32]
  wire  _T_11; // @[LZD.scala 39:14]
  wire  _T_12; // @[LZD.scala 39:21]
  wire  _T_13; // @[LZD.scala 39:30]
  wire  _T_14; // @[LZD.scala 39:27]
  wire  _T_15; // @[LZD.scala 39:25]
  wire [1:0] _T_16; // @[Cat.scala 29:58]
  wire [1:0] _T_17; // @[LZD.scala 44:32]
  wire  _T_18; // @[LZD.scala 39:14]
  wire  _T_19; // @[LZD.scala 39:21]
  wire  _T_20; // @[LZD.scala 39:30]
  wire  _T_21; // @[LZD.scala 39:27]
  wire  _T_22; // @[LZD.scala 39:25]
  wire [1:0] _T_23; // @[Cat.scala 29:58]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[Shift.scala 12:21]
  wire  _T_26; // @[LZD.scala 49:16]
  wire  _T_27; // @[LZD.scala 49:27]
  wire  _T_28; // @[LZD.scala 49:25]
  wire  _T_29; // @[LZD.scala 49:47]
  wire  _T_30; // @[LZD.scala 49:59]
  wire  _T_31; // @[LZD.scala 49:35]
  wire [2:0] _T_33; // @[Cat.scala 29:58]
  wire [3:0] _T_34; // @[LZD.scala 44:32]
  wire [1:0] _T_35; // @[LZD.scala 43:32]
  wire  _T_36; // @[LZD.scala 39:14]
  wire  _T_37; // @[LZD.scala 39:21]
  wire  _T_38; // @[LZD.scala 39:30]
  wire  _T_39; // @[LZD.scala 39:27]
  wire  _T_40; // @[LZD.scala 39:25]
  wire [1:0] _T_41; // @[Cat.scala 29:58]
  wire [1:0] _T_42; // @[LZD.scala 44:32]
  wire  _T_43; // @[LZD.scala 39:14]
  wire  _T_44; // @[LZD.scala 39:21]
  wire  _T_45; // @[LZD.scala 39:30]
  wire  _T_46; // @[LZD.scala 39:27]
  wire  _T_47; // @[LZD.scala 39:25]
  wire [1:0] _T_48; // @[Cat.scala 29:58]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[Shift.scala 12:21]
  wire  _T_51; // @[LZD.scala 49:16]
  wire  _T_52; // @[LZD.scala 49:27]
  wire  _T_53; // @[LZD.scala 49:25]
  wire  _T_54; // @[LZD.scala 49:47]
  wire  _T_55; // @[LZD.scala 49:59]
  wire  _T_56; // @[LZD.scala 49:35]
  wire [2:0] _T_58; // @[Cat.scala 29:58]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[LZD.scala 49:16]
  wire  _T_62; // @[LZD.scala 49:27]
  wire  _T_63; // @[LZD.scala 49:25]
  wire [1:0] _T_64; // @[LZD.scala 49:47]
  wire [1:0] _T_65; // @[LZD.scala 49:59]
  wire [1:0] _T_66; // @[LZD.scala 49:35]
  wire [3:0] _T_68; // @[Cat.scala 29:58]
  wire [7:0] _T_69; // @[LZD.scala 44:32]
  wire [3:0] _T_70; // @[LZD.scala 43:32]
  wire [1:0] _T_71; // @[LZD.scala 43:32]
  wire  _T_72; // @[LZD.scala 39:14]
  wire  _T_73; // @[LZD.scala 39:21]
  wire  _T_74; // @[LZD.scala 39:30]
  wire  _T_75; // @[LZD.scala 39:27]
  wire  _T_76; // @[LZD.scala 39:25]
  wire [1:0] _T_77; // @[Cat.scala 29:58]
  wire [1:0] _T_78; // @[LZD.scala 44:32]
  wire  _T_79; // @[LZD.scala 39:14]
  wire  _T_80; // @[LZD.scala 39:21]
  wire  _T_81; // @[LZD.scala 39:30]
  wire  _T_82; // @[LZD.scala 39:27]
  wire  _T_83; // @[LZD.scala 39:25]
  wire [1:0] _T_84; // @[Cat.scala 29:58]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[Shift.scala 12:21]
  wire  _T_87; // @[LZD.scala 49:16]
  wire  _T_88; // @[LZD.scala 49:27]
  wire  _T_89; // @[LZD.scala 49:25]
  wire  _T_90; // @[LZD.scala 49:47]
  wire  _T_91; // @[LZD.scala 49:59]
  wire  _T_92; // @[LZD.scala 49:35]
  wire [2:0] _T_94; // @[Cat.scala 29:58]
  wire [3:0] _T_95; // @[LZD.scala 44:32]
  wire [1:0] _T_96; // @[LZD.scala 43:32]
  wire  _T_97; // @[LZD.scala 39:14]
  wire  _T_98; // @[LZD.scala 39:21]
  wire  _T_99; // @[LZD.scala 39:30]
  wire  _T_100; // @[LZD.scala 39:27]
  wire  _T_101; // @[LZD.scala 39:25]
  wire [1:0] _T_102; // @[Cat.scala 29:58]
  wire [1:0] _T_103; // @[LZD.scala 44:32]
  wire  _T_104; // @[LZD.scala 39:14]
  wire  _T_105; // @[LZD.scala 39:21]
  wire  _T_106; // @[LZD.scala 39:30]
  wire  _T_107; // @[LZD.scala 39:27]
  wire  _T_108; // @[LZD.scala 39:25]
  wire [1:0] _T_109; // @[Cat.scala 29:58]
  wire  _T_110; // @[Shift.scala 12:21]
  wire  _T_111; // @[Shift.scala 12:21]
  wire  _T_112; // @[LZD.scala 49:16]
  wire  _T_113; // @[LZD.scala 49:27]
  wire  _T_114; // @[LZD.scala 49:25]
  wire  _T_115; // @[LZD.scala 49:47]
  wire  _T_116; // @[LZD.scala 49:59]
  wire  _T_117; // @[LZD.scala 49:35]
  wire [2:0] _T_119; // @[Cat.scala 29:58]
  wire  _T_120; // @[Shift.scala 12:21]
  wire  _T_121; // @[Shift.scala 12:21]
  wire  _T_122; // @[LZD.scala 49:16]
  wire  _T_123; // @[LZD.scala 49:27]
  wire  _T_124; // @[LZD.scala 49:25]
  wire [1:0] _T_125; // @[LZD.scala 49:47]
  wire [1:0] _T_126; // @[LZD.scala 49:59]
  wire [1:0] _T_127; // @[LZD.scala 49:35]
  wire [3:0] _T_129; // @[Cat.scala 29:58]
  wire  _T_130; // @[Shift.scala 12:21]
  wire  _T_131; // @[Shift.scala 12:21]
  wire  _T_132; // @[LZD.scala 49:16]
  wire  _T_133; // @[LZD.scala 49:27]
  wire  _T_134; // @[LZD.scala 49:25]
  wire [2:0] _T_135; // @[LZD.scala 49:47]
  wire [2:0] _T_136; // @[LZD.scala 49:59]
  wire [2:0] _T_137; // @[LZD.scala 49:35]
  wire [4:0] _T_139; // @[Cat.scala 29:58]
  wire [10:0] _T_140; // @[LZD.scala 44:32]
  wire [7:0] _T_141; // @[LZD.scala 43:32]
  wire [3:0] _T_142; // @[LZD.scala 43:32]
  wire [1:0] _T_143; // @[LZD.scala 43:32]
  wire  _T_144; // @[LZD.scala 39:14]
  wire  _T_145; // @[LZD.scala 39:21]
  wire  _T_146; // @[LZD.scala 39:30]
  wire  _T_147; // @[LZD.scala 39:27]
  wire  _T_148; // @[LZD.scala 39:25]
  wire [1:0] _T_149; // @[Cat.scala 29:58]
  wire [1:0] _T_150; // @[LZD.scala 44:32]
  wire  _T_151; // @[LZD.scala 39:14]
  wire  _T_152; // @[LZD.scala 39:21]
  wire  _T_153; // @[LZD.scala 39:30]
  wire  _T_154; // @[LZD.scala 39:27]
  wire  _T_155; // @[LZD.scala 39:25]
  wire [1:0] _T_156; // @[Cat.scala 29:58]
  wire  _T_157; // @[Shift.scala 12:21]
  wire  _T_158; // @[Shift.scala 12:21]
  wire  _T_159; // @[LZD.scala 49:16]
  wire  _T_160; // @[LZD.scala 49:27]
  wire  _T_161; // @[LZD.scala 49:25]
  wire  _T_162; // @[LZD.scala 49:47]
  wire  _T_163; // @[LZD.scala 49:59]
  wire  _T_164; // @[LZD.scala 49:35]
  wire [2:0] _T_166; // @[Cat.scala 29:58]
  wire [3:0] _T_167; // @[LZD.scala 44:32]
  wire [1:0] _T_168; // @[LZD.scala 43:32]
  wire  _T_169; // @[LZD.scala 39:14]
  wire  _T_170; // @[LZD.scala 39:21]
  wire  _T_171; // @[LZD.scala 39:30]
  wire  _T_172; // @[LZD.scala 39:27]
  wire  _T_173; // @[LZD.scala 39:25]
  wire [1:0] _T_174; // @[Cat.scala 29:58]
  wire [1:0] _T_175; // @[LZD.scala 44:32]
  wire  _T_176; // @[LZD.scala 39:14]
  wire  _T_177; // @[LZD.scala 39:21]
  wire  _T_178; // @[LZD.scala 39:30]
  wire  _T_179; // @[LZD.scala 39:27]
  wire  _T_180; // @[LZD.scala 39:25]
  wire [1:0] _T_181; // @[Cat.scala 29:58]
  wire  _T_182; // @[Shift.scala 12:21]
  wire  _T_183; // @[Shift.scala 12:21]
  wire  _T_184; // @[LZD.scala 49:16]
  wire  _T_185; // @[LZD.scala 49:27]
  wire  _T_186; // @[LZD.scala 49:25]
  wire  _T_187; // @[LZD.scala 49:47]
  wire  _T_188; // @[LZD.scala 49:59]
  wire  _T_189; // @[LZD.scala 49:35]
  wire [2:0] _T_191; // @[Cat.scala 29:58]
  wire  _T_192; // @[Shift.scala 12:21]
  wire  _T_193; // @[Shift.scala 12:21]
  wire  _T_194; // @[LZD.scala 49:16]
  wire  _T_195; // @[LZD.scala 49:27]
  wire  _T_196; // @[LZD.scala 49:25]
  wire [1:0] _T_197; // @[LZD.scala 49:47]
  wire [1:0] _T_198; // @[LZD.scala 49:59]
  wire [1:0] _T_199; // @[LZD.scala 49:35]
  wire [3:0] _T_201; // @[Cat.scala 29:58]
  wire [2:0] _T_202; // @[LZD.scala 44:32]
  wire [1:0] _T_203; // @[LZD.scala 43:32]
  wire  _T_204; // @[LZD.scala 39:14]
  wire  _T_205; // @[LZD.scala 39:21]
  wire  _T_206; // @[LZD.scala 39:30]
  wire  _T_207; // @[LZD.scala 39:27]
  wire  _T_208; // @[LZD.scala 39:25]
  wire [1:0] _T_209; // @[Cat.scala 29:58]
  wire  _T_210; // @[LZD.scala 44:32]
  wire  _T_212; // @[Shift.scala 12:21]
  wire  _T_214; // @[LZD.scala 55:32]
  wire  _T_215; // @[LZD.scala 55:20]
  wire  _T_217; // @[Shift.scala 12:21]
  wire [2:0] _T_219; // @[Cat.scala 29:58]
  wire [2:0] _T_220; // @[LZD.scala 55:32]
  wire [2:0] _T_221; // @[LZD.scala 55:20]
  wire [3:0] _T_222; // @[Cat.scala 29:58]
  wire  _T_223; // @[Shift.scala 12:21]
  wire [3:0] _T_225; // @[LZD.scala 55:32]
  wire [3:0] _T_226; // @[LZD.scala 55:20]
  wire [4:0] _T_227; // @[Cat.scala 29:58]
  wire [4:0] _T_228; // @[convert.scala 21:22]
  wire [25:0] _T_229; // @[convert.scala 22:36]
  wire  _T_230; // @[Shift.scala 16:24]
  wire  _T_232; // @[Shift.scala 12:21]
  wire [9:0] _T_233; // @[Shift.scala 64:52]
  wire [25:0] _T_235; // @[Cat.scala 29:58]
  wire [25:0] _T_236; // @[Shift.scala 64:27]
  wire [3:0] _T_237; // @[Shift.scala 66:70]
  wire  _T_238; // @[Shift.scala 12:21]
  wire [17:0] _T_239; // @[Shift.scala 64:52]
  wire [25:0] _T_241; // @[Cat.scala 29:58]
  wire [25:0] _T_242; // @[Shift.scala 64:27]
  wire [2:0] _T_243; // @[Shift.scala 66:70]
  wire  _T_244; // @[Shift.scala 12:21]
  wire [21:0] _T_245; // @[Shift.scala 64:52]
  wire [25:0] _T_247; // @[Cat.scala 29:58]
  wire [25:0] _T_248; // @[Shift.scala 64:27]
  wire [1:0] _T_249; // @[Shift.scala 66:70]
  wire  _T_250; // @[Shift.scala 12:21]
  wire [23:0] _T_251; // @[Shift.scala 64:52]
  wire [25:0] _T_253; // @[Cat.scala 29:58]
  wire [25:0] _T_254; // @[Shift.scala 64:27]
  wire  _T_255; // @[Shift.scala 66:70]
  wire [24:0] _T_257; // @[Shift.scala 64:52]
  wire [25:0] _T_258; // @[Cat.scala 29:58]
  wire [25:0] _T_259; // @[Shift.scala 64:27]
  wire [25:0] _T_260; // @[Shift.scala 16:10]
  wire [2:0] _T_261; // @[convert.scala 23:34]
  wire [22:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_263; // @[convert.scala 25:26]
  wire [4:0] _T_265; // @[convert.scala 25:42]
  wire [2:0] _T_268; // @[convert.scala 26:67]
  wire [2:0] _T_269; // @[convert.scala 26:51]
  wire [8:0] _T_270; // @[Cat.scala 29:58]
  wire [27:0] _T_272; // @[convert.scala 29:56]
  wire  _T_273; // @[convert.scala 29:60]
  wire  _T_274; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_277; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [8:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_286; // @[convert.scala 18:24]
  wire  _T_287; // @[convert.scala 18:40]
  wire  _T_288; // @[convert.scala 18:36]
  wire [26:0] _T_289; // @[convert.scala 19:24]
  wire [26:0] _T_290; // @[convert.scala 19:43]
  wire [26:0] _T_291; // @[convert.scala 19:39]
  wire [15:0] _T_292; // @[LZD.scala 43:32]
  wire [7:0] _T_293; // @[LZD.scala 43:32]
  wire [3:0] _T_294; // @[LZD.scala 43:32]
  wire [1:0] _T_295; // @[LZD.scala 43:32]
  wire  _T_296; // @[LZD.scala 39:14]
  wire  _T_297; // @[LZD.scala 39:21]
  wire  _T_298; // @[LZD.scala 39:30]
  wire  _T_299; // @[LZD.scala 39:27]
  wire  _T_300; // @[LZD.scala 39:25]
  wire [1:0] _T_301; // @[Cat.scala 29:58]
  wire [1:0] _T_302; // @[LZD.scala 44:32]
  wire  _T_303; // @[LZD.scala 39:14]
  wire  _T_304; // @[LZD.scala 39:21]
  wire  _T_305; // @[LZD.scala 39:30]
  wire  _T_306; // @[LZD.scala 39:27]
  wire  _T_307; // @[LZD.scala 39:25]
  wire [1:0] _T_308; // @[Cat.scala 29:58]
  wire  _T_309; // @[Shift.scala 12:21]
  wire  _T_310; // @[Shift.scala 12:21]
  wire  _T_311; // @[LZD.scala 49:16]
  wire  _T_312; // @[LZD.scala 49:27]
  wire  _T_313; // @[LZD.scala 49:25]
  wire  _T_314; // @[LZD.scala 49:47]
  wire  _T_315; // @[LZD.scala 49:59]
  wire  _T_316; // @[LZD.scala 49:35]
  wire [2:0] _T_318; // @[Cat.scala 29:58]
  wire [3:0] _T_319; // @[LZD.scala 44:32]
  wire [1:0] _T_320; // @[LZD.scala 43:32]
  wire  _T_321; // @[LZD.scala 39:14]
  wire  _T_322; // @[LZD.scala 39:21]
  wire  _T_323; // @[LZD.scala 39:30]
  wire  _T_324; // @[LZD.scala 39:27]
  wire  _T_325; // @[LZD.scala 39:25]
  wire [1:0] _T_326; // @[Cat.scala 29:58]
  wire [1:0] _T_327; // @[LZD.scala 44:32]
  wire  _T_328; // @[LZD.scala 39:14]
  wire  _T_329; // @[LZD.scala 39:21]
  wire  _T_330; // @[LZD.scala 39:30]
  wire  _T_331; // @[LZD.scala 39:27]
  wire  _T_332; // @[LZD.scala 39:25]
  wire [1:0] _T_333; // @[Cat.scala 29:58]
  wire  _T_334; // @[Shift.scala 12:21]
  wire  _T_335; // @[Shift.scala 12:21]
  wire  _T_336; // @[LZD.scala 49:16]
  wire  _T_337; // @[LZD.scala 49:27]
  wire  _T_338; // @[LZD.scala 49:25]
  wire  _T_339; // @[LZD.scala 49:47]
  wire  _T_340; // @[LZD.scala 49:59]
  wire  _T_341; // @[LZD.scala 49:35]
  wire [2:0] _T_343; // @[Cat.scala 29:58]
  wire  _T_344; // @[Shift.scala 12:21]
  wire  _T_345; // @[Shift.scala 12:21]
  wire  _T_346; // @[LZD.scala 49:16]
  wire  _T_347; // @[LZD.scala 49:27]
  wire  _T_348; // @[LZD.scala 49:25]
  wire [1:0] _T_349; // @[LZD.scala 49:47]
  wire [1:0] _T_350; // @[LZD.scala 49:59]
  wire [1:0] _T_351; // @[LZD.scala 49:35]
  wire [3:0] _T_353; // @[Cat.scala 29:58]
  wire [7:0] _T_354; // @[LZD.scala 44:32]
  wire [3:0] _T_355; // @[LZD.scala 43:32]
  wire [1:0] _T_356; // @[LZD.scala 43:32]
  wire  _T_357; // @[LZD.scala 39:14]
  wire  _T_358; // @[LZD.scala 39:21]
  wire  _T_359; // @[LZD.scala 39:30]
  wire  _T_360; // @[LZD.scala 39:27]
  wire  _T_361; // @[LZD.scala 39:25]
  wire [1:0] _T_362; // @[Cat.scala 29:58]
  wire [1:0] _T_363; // @[LZD.scala 44:32]
  wire  _T_364; // @[LZD.scala 39:14]
  wire  _T_365; // @[LZD.scala 39:21]
  wire  _T_366; // @[LZD.scala 39:30]
  wire  _T_367; // @[LZD.scala 39:27]
  wire  _T_368; // @[LZD.scala 39:25]
  wire [1:0] _T_369; // @[Cat.scala 29:58]
  wire  _T_370; // @[Shift.scala 12:21]
  wire  _T_371; // @[Shift.scala 12:21]
  wire  _T_372; // @[LZD.scala 49:16]
  wire  _T_373; // @[LZD.scala 49:27]
  wire  _T_374; // @[LZD.scala 49:25]
  wire  _T_375; // @[LZD.scala 49:47]
  wire  _T_376; // @[LZD.scala 49:59]
  wire  _T_377; // @[LZD.scala 49:35]
  wire [2:0] _T_379; // @[Cat.scala 29:58]
  wire [3:0] _T_380; // @[LZD.scala 44:32]
  wire [1:0] _T_381; // @[LZD.scala 43:32]
  wire  _T_382; // @[LZD.scala 39:14]
  wire  _T_383; // @[LZD.scala 39:21]
  wire  _T_384; // @[LZD.scala 39:30]
  wire  _T_385; // @[LZD.scala 39:27]
  wire  _T_386; // @[LZD.scala 39:25]
  wire [1:0] _T_387; // @[Cat.scala 29:58]
  wire [1:0] _T_388; // @[LZD.scala 44:32]
  wire  _T_389; // @[LZD.scala 39:14]
  wire  _T_390; // @[LZD.scala 39:21]
  wire  _T_391; // @[LZD.scala 39:30]
  wire  _T_392; // @[LZD.scala 39:27]
  wire  _T_393; // @[LZD.scala 39:25]
  wire [1:0] _T_394; // @[Cat.scala 29:58]
  wire  _T_395; // @[Shift.scala 12:21]
  wire  _T_396; // @[Shift.scala 12:21]
  wire  _T_397; // @[LZD.scala 49:16]
  wire  _T_398; // @[LZD.scala 49:27]
  wire  _T_399; // @[LZD.scala 49:25]
  wire  _T_400; // @[LZD.scala 49:47]
  wire  _T_401; // @[LZD.scala 49:59]
  wire  _T_402; // @[LZD.scala 49:35]
  wire [2:0] _T_404; // @[Cat.scala 29:58]
  wire  _T_405; // @[Shift.scala 12:21]
  wire  _T_406; // @[Shift.scala 12:21]
  wire  _T_407; // @[LZD.scala 49:16]
  wire  _T_408; // @[LZD.scala 49:27]
  wire  _T_409; // @[LZD.scala 49:25]
  wire [1:0] _T_410; // @[LZD.scala 49:47]
  wire [1:0] _T_411; // @[LZD.scala 49:59]
  wire [1:0] _T_412; // @[LZD.scala 49:35]
  wire [3:0] _T_414; // @[Cat.scala 29:58]
  wire  _T_415; // @[Shift.scala 12:21]
  wire  _T_416; // @[Shift.scala 12:21]
  wire  _T_417; // @[LZD.scala 49:16]
  wire  _T_418; // @[LZD.scala 49:27]
  wire  _T_419; // @[LZD.scala 49:25]
  wire [2:0] _T_420; // @[LZD.scala 49:47]
  wire [2:0] _T_421; // @[LZD.scala 49:59]
  wire [2:0] _T_422; // @[LZD.scala 49:35]
  wire [4:0] _T_424; // @[Cat.scala 29:58]
  wire [10:0] _T_425; // @[LZD.scala 44:32]
  wire [7:0] _T_426; // @[LZD.scala 43:32]
  wire [3:0] _T_427; // @[LZD.scala 43:32]
  wire [1:0] _T_428; // @[LZD.scala 43:32]
  wire  _T_429; // @[LZD.scala 39:14]
  wire  _T_430; // @[LZD.scala 39:21]
  wire  _T_431; // @[LZD.scala 39:30]
  wire  _T_432; // @[LZD.scala 39:27]
  wire  _T_433; // @[LZD.scala 39:25]
  wire [1:0] _T_434; // @[Cat.scala 29:58]
  wire [1:0] _T_435; // @[LZD.scala 44:32]
  wire  _T_436; // @[LZD.scala 39:14]
  wire  _T_437; // @[LZD.scala 39:21]
  wire  _T_438; // @[LZD.scala 39:30]
  wire  _T_439; // @[LZD.scala 39:27]
  wire  _T_440; // @[LZD.scala 39:25]
  wire [1:0] _T_441; // @[Cat.scala 29:58]
  wire  _T_442; // @[Shift.scala 12:21]
  wire  _T_443; // @[Shift.scala 12:21]
  wire  _T_444; // @[LZD.scala 49:16]
  wire  _T_445; // @[LZD.scala 49:27]
  wire  _T_446; // @[LZD.scala 49:25]
  wire  _T_447; // @[LZD.scala 49:47]
  wire  _T_448; // @[LZD.scala 49:59]
  wire  _T_449; // @[LZD.scala 49:35]
  wire [2:0] _T_451; // @[Cat.scala 29:58]
  wire [3:0] _T_452; // @[LZD.scala 44:32]
  wire [1:0] _T_453; // @[LZD.scala 43:32]
  wire  _T_454; // @[LZD.scala 39:14]
  wire  _T_455; // @[LZD.scala 39:21]
  wire  _T_456; // @[LZD.scala 39:30]
  wire  _T_457; // @[LZD.scala 39:27]
  wire  _T_458; // @[LZD.scala 39:25]
  wire [1:0] _T_459; // @[Cat.scala 29:58]
  wire [1:0] _T_460; // @[LZD.scala 44:32]
  wire  _T_461; // @[LZD.scala 39:14]
  wire  _T_462; // @[LZD.scala 39:21]
  wire  _T_463; // @[LZD.scala 39:30]
  wire  _T_464; // @[LZD.scala 39:27]
  wire  _T_465; // @[LZD.scala 39:25]
  wire [1:0] _T_466; // @[Cat.scala 29:58]
  wire  _T_467; // @[Shift.scala 12:21]
  wire  _T_468; // @[Shift.scala 12:21]
  wire  _T_469; // @[LZD.scala 49:16]
  wire  _T_470; // @[LZD.scala 49:27]
  wire  _T_471; // @[LZD.scala 49:25]
  wire  _T_472; // @[LZD.scala 49:47]
  wire  _T_473; // @[LZD.scala 49:59]
  wire  _T_474; // @[LZD.scala 49:35]
  wire [2:0] _T_476; // @[Cat.scala 29:58]
  wire  _T_477; // @[Shift.scala 12:21]
  wire  _T_478; // @[Shift.scala 12:21]
  wire  _T_479; // @[LZD.scala 49:16]
  wire  _T_480; // @[LZD.scala 49:27]
  wire  _T_481; // @[LZD.scala 49:25]
  wire [1:0] _T_482; // @[LZD.scala 49:47]
  wire [1:0] _T_483; // @[LZD.scala 49:59]
  wire [1:0] _T_484; // @[LZD.scala 49:35]
  wire [3:0] _T_486; // @[Cat.scala 29:58]
  wire [2:0] _T_487; // @[LZD.scala 44:32]
  wire [1:0] _T_488; // @[LZD.scala 43:32]
  wire  _T_489; // @[LZD.scala 39:14]
  wire  _T_490; // @[LZD.scala 39:21]
  wire  _T_491; // @[LZD.scala 39:30]
  wire  _T_492; // @[LZD.scala 39:27]
  wire  _T_493; // @[LZD.scala 39:25]
  wire [1:0] _T_494; // @[Cat.scala 29:58]
  wire  _T_495; // @[LZD.scala 44:32]
  wire  _T_497; // @[Shift.scala 12:21]
  wire  _T_499; // @[LZD.scala 55:32]
  wire  _T_500; // @[LZD.scala 55:20]
  wire  _T_502; // @[Shift.scala 12:21]
  wire [2:0] _T_504; // @[Cat.scala 29:58]
  wire [2:0] _T_505; // @[LZD.scala 55:32]
  wire [2:0] _T_506; // @[LZD.scala 55:20]
  wire [3:0] _T_507; // @[Cat.scala 29:58]
  wire  _T_508; // @[Shift.scala 12:21]
  wire [3:0] _T_510; // @[LZD.scala 55:32]
  wire [3:0] _T_511; // @[LZD.scala 55:20]
  wire [4:0] _T_512; // @[Cat.scala 29:58]
  wire [4:0] _T_513; // @[convert.scala 21:22]
  wire [25:0] _T_514; // @[convert.scala 22:36]
  wire  _T_515; // @[Shift.scala 16:24]
  wire  _T_517; // @[Shift.scala 12:21]
  wire [9:0] _T_518; // @[Shift.scala 64:52]
  wire [25:0] _T_520; // @[Cat.scala 29:58]
  wire [25:0] _T_521; // @[Shift.scala 64:27]
  wire [3:0] _T_522; // @[Shift.scala 66:70]
  wire  _T_523; // @[Shift.scala 12:21]
  wire [17:0] _T_524; // @[Shift.scala 64:52]
  wire [25:0] _T_526; // @[Cat.scala 29:58]
  wire [25:0] _T_527; // @[Shift.scala 64:27]
  wire [2:0] _T_528; // @[Shift.scala 66:70]
  wire  _T_529; // @[Shift.scala 12:21]
  wire [21:0] _T_530; // @[Shift.scala 64:52]
  wire [25:0] _T_532; // @[Cat.scala 29:58]
  wire [25:0] _T_533; // @[Shift.scala 64:27]
  wire [1:0] _T_534; // @[Shift.scala 66:70]
  wire  _T_535; // @[Shift.scala 12:21]
  wire [23:0] _T_536; // @[Shift.scala 64:52]
  wire [25:0] _T_538; // @[Cat.scala 29:58]
  wire [25:0] _T_539; // @[Shift.scala 64:27]
  wire  _T_540; // @[Shift.scala 66:70]
  wire [24:0] _T_542; // @[Shift.scala 64:52]
  wire [25:0] _T_543; // @[Cat.scala 29:58]
  wire [25:0] _T_544; // @[Shift.scala 64:27]
  wire [25:0] _T_545; // @[Shift.scala 16:10]
  wire [2:0] _T_546; // @[convert.scala 23:34]
  wire [22:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_548; // @[convert.scala 25:26]
  wire [4:0] _T_550; // @[convert.scala 25:42]
  wire [2:0] _T_553; // @[convert.scala 26:67]
  wire [2:0] _T_554; // @[convert.scala 26:51]
  wire [8:0] _T_555; // @[Cat.scala 29:58]
  wire [27:0] _T_557; // @[convert.scala 29:56]
  wire  _T_558; // @[convert.scala 29:60]
  wire  _T_559; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_562; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [8:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[PositAdder.scala 24:32]
  wire  greaterSign; // @[PositAdder.scala 25:24]
  wire  smallerSign; // @[PositAdder.scala 26:24]
  wire [8:0] greaterExp; // @[PositAdder.scala 27:24]
  wire [8:0] smallerExp; // @[PositAdder.scala 28:24]
  wire [22:0] greaterFrac; // @[PositAdder.scala 29:24]
  wire [22:0] smallerFrac; // @[PositAdder.scala 30:24]
  wire [8:0] _T_571; // @[PositAdder.scala 31:32]
  wire [8:0] scale_diff; // @[PositAdder.scala 31:32]
  wire  _T_572; // @[PositAdder.scala 32:38]
  wire [24:0] greaterSig; // @[Cat.scala 29:58]
  wire  _T_574; // @[PositAdder.scala 33:38]
  wire [27:0] _T_577; // @[Cat.scala 29:58]
  wire [8:0] _T_578; // @[PositAdder.scala 34:68]
  wire  _T_579; // @[Shift.scala 39:24]
  wire [4:0] _T_580; // @[Shift.scala 40:44]
  wire [11:0] _T_581; // @[Shift.scala 90:30]
  wire [15:0] _T_582; // @[Shift.scala 90:48]
  wire  _T_583; // @[Shift.scala 90:57]
  wire [11:0] _GEN_0; // @[Shift.scala 90:39]
  wire [11:0] _T_584; // @[Shift.scala 90:39]
  wire  _T_585; // @[Shift.scala 12:21]
  wire  _T_586; // @[Shift.scala 12:21]
  wire [15:0] _T_588; // @[Bitwise.scala 71:12]
  wire [27:0] _T_589; // @[Cat.scala 29:58]
  wire [27:0] _T_590; // @[Shift.scala 91:22]
  wire [3:0] _T_591; // @[Shift.scala 92:77]
  wire [19:0] _T_592; // @[Shift.scala 90:30]
  wire [7:0] _T_593; // @[Shift.scala 90:48]
  wire  _T_594; // @[Shift.scala 90:57]
  wire [19:0] _GEN_1; // @[Shift.scala 90:39]
  wire [19:0] _T_595; // @[Shift.scala 90:39]
  wire  _T_596; // @[Shift.scala 12:21]
  wire  _T_597; // @[Shift.scala 12:21]
  wire [7:0] _T_599; // @[Bitwise.scala 71:12]
  wire [27:0] _T_600; // @[Cat.scala 29:58]
  wire [27:0] _T_601; // @[Shift.scala 91:22]
  wire [2:0] _T_602; // @[Shift.scala 92:77]
  wire [23:0] _T_603; // @[Shift.scala 90:30]
  wire [3:0] _T_604; // @[Shift.scala 90:48]
  wire  _T_605; // @[Shift.scala 90:57]
  wire [23:0] _GEN_2; // @[Shift.scala 90:39]
  wire [23:0] _T_606; // @[Shift.scala 90:39]
  wire  _T_607; // @[Shift.scala 12:21]
  wire  _T_608; // @[Shift.scala 12:21]
  wire [3:0] _T_610; // @[Bitwise.scala 71:12]
  wire [27:0] _T_611; // @[Cat.scala 29:58]
  wire [27:0] _T_612; // @[Shift.scala 91:22]
  wire [1:0] _T_613; // @[Shift.scala 92:77]
  wire [25:0] _T_614; // @[Shift.scala 90:30]
  wire [1:0] _T_615; // @[Shift.scala 90:48]
  wire  _T_616; // @[Shift.scala 90:57]
  wire [25:0] _GEN_3; // @[Shift.scala 90:39]
  wire [25:0] _T_617; // @[Shift.scala 90:39]
  wire  _T_618; // @[Shift.scala 12:21]
  wire  _T_619; // @[Shift.scala 12:21]
  wire [1:0] _T_621; // @[Bitwise.scala 71:12]
  wire [27:0] _T_622; // @[Cat.scala 29:58]
  wire [27:0] _T_623; // @[Shift.scala 91:22]
  wire  _T_624; // @[Shift.scala 92:77]
  wire [26:0] _T_625; // @[Shift.scala 90:30]
  wire  _T_626; // @[Shift.scala 90:48]
  wire [26:0] _GEN_4; // @[Shift.scala 90:39]
  wire [26:0] _T_628; // @[Shift.scala 90:39]
  wire  _T_630; // @[Shift.scala 12:21]
  wire [27:0] _T_631; // @[Cat.scala 29:58]
  wire [27:0] _T_632; // @[Shift.scala 91:22]
  wire [27:0] _T_635; // @[Bitwise.scala 71:12]
  wire [27:0] smallerSig; // @[Shift.scala 39:10]
  wire [24:0] _T_636; // @[PositAdder.scala 35:45]
  wire [25:0] rawSumSig; // @[PositAdder.scala 35:32]
  wire  _T_637; // @[PositAdder.scala 36:31]
  wire  _T_638; // @[PositAdder.scala 36:59]
  wire  sumSign; // @[PositAdder.scala 36:43]
  wire [24:0] _T_639; // @[PositAdder.scala 37:48]
  wire [2:0] _T_640; // @[PositAdder.scala 37:63]
  wire [28:0] signSumSig; // @[Cat.scala 29:58]
  wire [27:0] _T_642; // @[PositAdder.scala 39:31]
  wire [27:0] _T_643; // @[PositAdder.scala 39:66]
  wire [27:0] sumXor; // @[PositAdder.scala 39:49]
  wire [15:0] _T_644; // @[LZD.scala 43:32]
  wire [7:0] _T_645; // @[LZD.scala 43:32]
  wire [3:0] _T_646; // @[LZD.scala 43:32]
  wire [1:0] _T_647; // @[LZD.scala 43:32]
  wire  _T_648; // @[LZD.scala 39:14]
  wire  _T_649; // @[LZD.scala 39:21]
  wire  _T_650; // @[LZD.scala 39:30]
  wire  _T_651; // @[LZD.scala 39:27]
  wire  _T_652; // @[LZD.scala 39:25]
  wire [1:0] _T_653; // @[Cat.scala 29:58]
  wire [1:0] _T_654; // @[LZD.scala 44:32]
  wire  _T_655; // @[LZD.scala 39:14]
  wire  _T_656; // @[LZD.scala 39:21]
  wire  _T_657; // @[LZD.scala 39:30]
  wire  _T_658; // @[LZD.scala 39:27]
  wire  _T_659; // @[LZD.scala 39:25]
  wire [1:0] _T_660; // @[Cat.scala 29:58]
  wire  _T_661; // @[Shift.scala 12:21]
  wire  _T_662; // @[Shift.scala 12:21]
  wire  _T_663; // @[LZD.scala 49:16]
  wire  _T_664; // @[LZD.scala 49:27]
  wire  _T_665; // @[LZD.scala 49:25]
  wire  _T_666; // @[LZD.scala 49:47]
  wire  _T_667; // @[LZD.scala 49:59]
  wire  _T_668; // @[LZD.scala 49:35]
  wire [2:0] _T_670; // @[Cat.scala 29:58]
  wire [3:0] _T_671; // @[LZD.scala 44:32]
  wire [1:0] _T_672; // @[LZD.scala 43:32]
  wire  _T_673; // @[LZD.scala 39:14]
  wire  _T_674; // @[LZD.scala 39:21]
  wire  _T_675; // @[LZD.scala 39:30]
  wire  _T_676; // @[LZD.scala 39:27]
  wire  _T_677; // @[LZD.scala 39:25]
  wire [1:0] _T_678; // @[Cat.scala 29:58]
  wire [1:0] _T_679; // @[LZD.scala 44:32]
  wire  _T_680; // @[LZD.scala 39:14]
  wire  _T_681; // @[LZD.scala 39:21]
  wire  _T_682; // @[LZD.scala 39:30]
  wire  _T_683; // @[LZD.scala 39:27]
  wire  _T_684; // @[LZD.scala 39:25]
  wire [1:0] _T_685; // @[Cat.scala 29:58]
  wire  _T_686; // @[Shift.scala 12:21]
  wire  _T_687; // @[Shift.scala 12:21]
  wire  _T_688; // @[LZD.scala 49:16]
  wire  _T_689; // @[LZD.scala 49:27]
  wire  _T_690; // @[LZD.scala 49:25]
  wire  _T_691; // @[LZD.scala 49:47]
  wire  _T_692; // @[LZD.scala 49:59]
  wire  _T_693; // @[LZD.scala 49:35]
  wire [2:0] _T_695; // @[Cat.scala 29:58]
  wire  _T_696; // @[Shift.scala 12:21]
  wire  _T_697; // @[Shift.scala 12:21]
  wire  _T_698; // @[LZD.scala 49:16]
  wire  _T_699; // @[LZD.scala 49:27]
  wire  _T_700; // @[LZD.scala 49:25]
  wire [1:0] _T_701; // @[LZD.scala 49:47]
  wire [1:0] _T_702; // @[LZD.scala 49:59]
  wire [1:0] _T_703; // @[LZD.scala 49:35]
  wire [3:0] _T_705; // @[Cat.scala 29:58]
  wire [7:0] _T_706; // @[LZD.scala 44:32]
  wire [3:0] _T_707; // @[LZD.scala 43:32]
  wire [1:0] _T_708; // @[LZD.scala 43:32]
  wire  _T_709; // @[LZD.scala 39:14]
  wire  _T_710; // @[LZD.scala 39:21]
  wire  _T_711; // @[LZD.scala 39:30]
  wire  _T_712; // @[LZD.scala 39:27]
  wire  _T_713; // @[LZD.scala 39:25]
  wire [1:0] _T_714; // @[Cat.scala 29:58]
  wire [1:0] _T_715; // @[LZD.scala 44:32]
  wire  _T_716; // @[LZD.scala 39:14]
  wire  _T_717; // @[LZD.scala 39:21]
  wire  _T_718; // @[LZD.scala 39:30]
  wire  _T_719; // @[LZD.scala 39:27]
  wire  _T_720; // @[LZD.scala 39:25]
  wire [1:0] _T_721; // @[Cat.scala 29:58]
  wire  _T_722; // @[Shift.scala 12:21]
  wire  _T_723; // @[Shift.scala 12:21]
  wire  _T_724; // @[LZD.scala 49:16]
  wire  _T_725; // @[LZD.scala 49:27]
  wire  _T_726; // @[LZD.scala 49:25]
  wire  _T_727; // @[LZD.scala 49:47]
  wire  _T_728; // @[LZD.scala 49:59]
  wire  _T_729; // @[LZD.scala 49:35]
  wire [2:0] _T_731; // @[Cat.scala 29:58]
  wire [3:0] _T_732; // @[LZD.scala 44:32]
  wire [1:0] _T_733; // @[LZD.scala 43:32]
  wire  _T_734; // @[LZD.scala 39:14]
  wire  _T_735; // @[LZD.scala 39:21]
  wire  _T_736; // @[LZD.scala 39:30]
  wire  _T_737; // @[LZD.scala 39:27]
  wire  _T_738; // @[LZD.scala 39:25]
  wire [1:0] _T_739; // @[Cat.scala 29:58]
  wire [1:0] _T_740; // @[LZD.scala 44:32]
  wire  _T_741; // @[LZD.scala 39:14]
  wire  _T_742; // @[LZD.scala 39:21]
  wire  _T_743; // @[LZD.scala 39:30]
  wire  _T_744; // @[LZD.scala 39:27]
  wire  _T_745; // @[LZD.scala 39:25]
  wire [1:0] _T_746; // @[Cat.scala 29:58]
  wire  _T_747; // @[Shift.scala 12:21]
  wire  _T_748; // @[Shift.scala 12:21]
  wire  _T_749; // @[LZD.scala 49:16]
  wire  _T_750; // @[LZD.scala 49:27]
  wire  _T_751; // @[LZD.scala 49:25]
  wire  _T_752; // @[LZD.scala 49:47]
  wire  _T_753; // @[LZD.scala 49:59]
  wire  _T_754; // @[LZD.scala 49:35]
  wire [2:0] _T_756; // @[Cat.scala 29:58]
  wire  _T_757; // @[Shift.scala 12:21]
  wire  _T_758; // @[Shift.scala 12:21]
  wire  _T_759; // @[LZD.scala 49:16]
  wire  _T_760; // @[LZD.scala 49:27]
  wire  _T_761; // @[LZD.scala 49:25]
  wire [1:0] _T_762; // @[LZD.scala 49:47]
  wire [1:0] _T_763; // @[LZD.scala 49:59]
  wire [1:0] _T_764; // @[LZD.scala 49:35]
  wire [3:0] _T_766; // @[Cat.scala 29:58]
  wire  _T_767; // @[Shift.scala 12:21]
  wire  _T_768; // @[Shift.scala 12:21]
  wire  _T_769; // @[LZD.scala 49:16]
  wire  _T_770; // @[LZD.scala 49:27]
  wire  _T_771; // @[LZD.scala 49:25]
  wire [2:0] _T_772; // @[LZD.scala 49:47]
  wire [2:0] _T_773; // @[LZD.scala 49:59]
  wire [2:0] _T_774; // @[LZD.scala 49:35]
  wire [4:0] _T_776; // @[Cat.scala 29:58]
  wire [11:0] _T_777; // @[LZD.scala 44:32]
  wire [7:0] _T_778; // @[LZD.scala 43:32]
  wire [3:0] _T_779; // @[LZD.scala 43:32]
  wire [1:0] _T_780; // @[LZD.scala 43:32]
  wire  _T_781; // @[LZD.scala 39:14]
  wire  _T_782; // @[LZD.scala 39:21]
  wire  _T_783; // @[LZD.scala 39:30]
  wire  _T_784; // @[LZD.scala 39:27]
  wire  _T_785; // @[LZD.scala 39:25]
  wire [1:0] _T_786; // @[Cat.scala 29:58]
  wire [1:0] _T_787; // @[LZD.scala 44:32]
  wire  _T_788; // @[LZD.scala 39:14]
  wire  _T_789; // @[LZD.scala 39:21]
  wire  _T_790; // @[LZD.scala 39:30]
  wire  _T_791; // @[LZD.scala 39:27]
  wire  _T_792; // @[LZD.scala 39:25]
  wire [1:0] _T_793; // @[Cat.scala 29:58]
  wire  _T_794; // @[Shift.scala 12:21]
  wire  _T_795; // @[Shift.scala 12:21]
  wire  _T_796; // @[LZD.scala 49:16]
  wire  _T_797; // @[LZD.scala 49:27]
  wire  _T_798; // @[LZD.scala 49:25]
  wire  _T_799; // @[LZD.scala 49:47]
  wire  _T_800; // @[LZD.scala 49:59]
  wire  _T_801; // @[LZD.scala 49:35]
  wire [2:0] _T_803; // @[Cat.scala 29:58]
  wire [3:0] _T_804; // @[LZD.scala 44:32]
  wire [1:0] _T_805; // @[LZD.scala 43:32]
  wire  _T_806; // @[LZD.scala 39:14]
  wire  _T_807; // @[LZD.scala 39:21]
  wire  _T_808; // @[LZD.scala 39:30]
  wire  _T_809; // @[LZD.scala 39:27]
  wire  _T_810; // @[LZD.scala 39:25]
  wire [1:0] _T_811; // @[Cat.scala 29:58]
  wire [1:0] _T_812; // @[LZD.scala 44:32]
  wire  _T_813; // @[LZD.scala 39:14]
  wire  _T_814; // @[LZD.scala 39:21]
  wire  _T_815; // @[LZD.scala 39:30]
  wire  _T_816; // @[LZD.scala 39:27]
  wire  _T_817; // @[LZD.scala 39:25]
  wire [1:0] _T_818; // @[Cat.scala 29:58]
  wire  _T_819; // @[Shift.scala 12:21]
  wire  _T_820; // @[Shift.scala 12:21]
  wire  _T_821; // @[LZD.scala 49:16]
  wire  _T_822; // @[LZD.scala 49:27]
  wire  _T_823; // @[LZD.scala 49:25]
  wire  _T_824; // @[LZD.scala 49:47]
  wire  _T_825; // @[LZD.scala 49:59]
  wire  _T_826; // @[LZD.scala 49:35]
  wire [2:0] _T_828; // @[Cat.scala 29:58]
  wire  _T_829; // @[Shift.scala 12:21]
  wire  _T_830; // @[Shift.scala 12:21]
  wire  _T_831; // @[LZD.scala 49:16]
  wire  _T_832; // @[LZD.scala 49:27]
  wire  _T_833; // @[LZD.scala 49:25]
  wire [1:0] _T_834; // @[LZD.scala 49:47]
  wire [1:0] _T_835; // @[LZD.scala 49:59]
  wire [1:0] _T_836; // @[LZD.scala 49:35]
  wire [3:0] _T_838; // @[Cat.scala 29:58]
  wire [3:0] _T_839; // @[LZD.scala 44:32]
  wire [1:0] _T_840; // @[LZD.scala 43:32]
  wire  _T_841; // @[LZD.scala 39:14]
  wire  _T_842; // @[LZD.scala 39:21]
  wire  _T_843; // @[LZD.scala 39:30]
  wire  _T_844; // @[LZD.scala 39:27]
  wire  _T_845; // @[LZD.scala 39:25]
  wire [1:0] _T_846; // @[Cat.scala 29:58]
  wire [1:0] _T_847; // @[LZD.scala 44:32]
  wire  _T_848; // @[LZD.scala 39:14]
  wire  _T_849; // @[LZD.scala 39:21]
  wire  _T_850; // @[LZD.scala 39:30]
  wire  _T_851; // @[LZD.scala 39:27]
  wire  _T_852; // @[LZD.scala 39:25]
  wire [1:0] _T_853; // @[Cat.scala 29:58]
  wire  _T_854; // @[Shift.scala 12:21]
  wire  _T_855; // @[Shift.scala 12:21]
  wire  _T_856; // @[LZD.scala 49:16]
  wire  _T_857; // @[LZD.scala 49:27]
  wire  _T_858; // @[LZD.scala 49:25]
  wire  _T_859; // @[LZD.scala 49:47]
  wire  _T_860; // @[LZD.scala 49:59]
  wire  _T_861; // @[LZD.scala 49:35]
  wire [2:0] _T_863; // @[Cat.scala 29:58]
  wire  _T_864; // @[Shift.scala 12:21]
  wire [2:0] _T_866; // @[LZD.scala 55:32]
  wire [2:0] _T_867; // @[LZD.scala 55:20]
  wire [3:0] _T_868; // @[Cat.scala 29:58]
  wire  _T_869; // @[Shift.scala 12:21]
  wire [3:0] _T_871; // @[LZD.scala 55:32]
  wire [3:0] _T_872; // @[LZD.scala 55:20]
  wire [4:0] sumLZD; // @[Cat.scala 29:58]
  wire [5:0] _T_873; // @[Cat.scala 29:58]
  wire [5:0] _T_874; // @[PositAdder.scala 41:38]
  wire [5:0] _T_876; // @[PositAdder.scala 41:45]
  wire [5:0] scaleBias; // @[PositAdder.scala 41:45]
  wire [8:0] _GEN_5; // @[PositAdder.scala 42:32]
  wire [9:0] sumScale; // @[PositAdder.scala 42:32]
  wire  overflow; // @[PositAdder.scala 43:30]
  wire [4:0] normalShift; // @[PositAdder.scala 44:22]
  wire [26:0] _T_877; // @[PositAdder.scala 45:36]
  wire  _T_878; // @[Shift.scala 16:24]
  wire  _T_880; // @[Shift.scala 12:21]
  wire [10:0] _T_881; // @[Shift.scala 64:52]
  wire [26:0] _T_883; // @[Cat.scala 29:58]
  wire [26:0] _T_884; // @[Shift.scala 64:27]
  wire [3:0] _T_885; // @[Shift.scala 66:70]
  wire  _T_886; // @[Shift.scala 12:21]
  wire [18:0] _T_887; // @[Shift.scala 64:52]
  wire [26:0] _T_889; // @[Cat.scala 29:58]
  wire [26:0] _T_890; // @[Shift.scala 64:27]
  wire [2:0] _T_891; // @[Shift.scala 66:70]
  wire  _T_892; // @[Shift.scala 12:21]
  wire [22:0] _T_893; // @[Shift.scala 64:52]
  wire [26:0] _T_895; // @[Cat.scala 29:58]
  wire [26:0] _T_896; // @[Shift.scala 64:27]
  wire [1:0] _T_897; // @[Shift.scala 66:70]
  wire  _T_898; // @[Shift.scala 12:21]
  wire [24:0] _T_899; // @[Shift.scala 64:52]
  wire [26:0] _T_901; // @[Cat.scala 29:58]
  wire [26:0] _T_902; // @[Shift.scala 64:27]
  wire  _T_903; // @[Shift.scala 66:70]
  wire [25:0] _T_905; // @[Shift.scala 64:52]
  wire [26:0] _T_906; // @[Cat.scala 29:58]
  wire [26:0] _T_907; // @[Shift.scala 64:27]
  wire [26:0] shiftSig; // @[Shift.scala 16:10]
  wire [9:0] _T_908; // @[PositAdder.scala 50:24]
  wire [22:0] decS_fraction; // @[PositAdder.scala 51:34]
  wire  decS_isNaR; // @[PositAdder.scala 52:32]
  wire  _T_911; // @[PositAdder.scala 53:33]
  wire  _T_912; // @[PositAdder.scala 53:21]
  wire  _T_913; // @[PositAdder.scala 53:52]
  wire  decS_isZero; // @[PositAdder.scala 53:37]
  wire [1:0] _T_915; // @[PositAdder.scala 54:33]
  wire  _T_916; // @[PositAdder.scala 54:49]
  wire  _T_917; // @[PositAdder.scala 54:63]
  wire  _T_918; // @[PositAdder.scala 54:53]
  wire [8:0] _GEN_6; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  wire [8:0] decS_scale; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  wire [2:0] _T_921; // @[convert.scala 46:61]
  wire [2:0] _T_922; // @[convert.scala 46:52]
  wire [2:0] _T_924; // @[convert.scala 46:42]
  wire [5:0] _T_925; // @[convert.scala 48:34]
  wire  _T_926; // @[convert.scala 49:36]
  wire [5:0] _T_928; // @[convert.scala 50:36]
  wire [5:0] _T_929; // @[convert.scala 50:36]
  wire [5:0] _T_930; // @[convert.scala 50:28]
  wire  _T_931; // @[convert.scala 51:31]
  wire  _T_932; // @[convert.scala 52:43]
  wire [30:0] _T_936; // @[Cat.scala 29:58]
  wire [5:0] _T_937; // @[Shift.scala 39:17]
  wire  _T_938; // @[Shift.scala 39:24]
  wire [4:0] _T_939; // @[Shift.scala 40:44]
  wire [14:0] _T_940; // @[Shift.scala 90:30]
  wire [15:0] _T_941; // @[Shift.scala 90:48]
  wire  _T_942; // @[Shift.scala 90:57]
  wire [14:0] _GEN_7; // @[Shift.scala 90:39]
  wire [14:0] _T_943; // @[Shift.scala 90:39]
  wire  _T_944; // @[Shift.scala 12:21]
  wire  _T_945; // @[Shift.scala 12:21]
  wire [15:0] _T_947; // @[Bitwise.scala 71:12]
  wire [30:0] _T_948; // @[Cat.scala 29:58]
  wire [30:0] _T_949; // @[Shift.scala 91:22]
  wire [3:0] _T_950; // @[Shift.scala 92:77]
  wire [22:0] _T_951; // @[Shift.scala 90:30]
  wire [7:0] _T_952; // @[Shift.scala 90:48]
  wire  _T_953; // @[Shift.scala 90:57]
  wire [22:0] _GEN_8; // @[Shift.scala 90:39]
  wire [22:0] _T_954; // @[Shift.scala 90:39]
  wire  _T_955; // @[Shift.scala 12:21]
  wire  _T_956; // @[Shift.scala 12:21]
  wire [7:0] _T_958; // @[Bitwise.scala 71:12]
  wire [30:0] _T_959; // @[Cat.scala 29:58]
  wire [30:0] _T_960; // @[Shift.scala 91:22]
  wire [2:0] _T_961; // @[Shift.scala 92:77]
  wire [26:0] _T_962; // @[Shift.scala 90:30]
  wire [3:0] _T_963; // @[Shift.scala 90:48]
  wire  _T_964; // @[Shift.scala 90:57]
  wire [26:0] _GEN_9; // @[Shift.scala 90:39]
  wire [26:0] _T_965; // @[Shift.scala 90:39]
  wire  _T_966; // @[Shift.scala 12:21]
  wire  _T_967; // @[Shift.scala 12:21]
  wire [3:0] _T_969; // @[Bitwise.scala 71:12]
  wire [30:0] _T_970; // @[Cat.scala 29:58]
  wire [30:0] _T_971; // @[Shift.scala 91:22]
  wire [1:0] _T_972; // @[Shift.scala 92:77]
  wire [28:0] _T_973; // @[Shift.scala 90:30]
  wire [1:0] _T_974; // @[Shift.scala 90:48]
  wire  _T_975; // @[Shift.scala 90:57]
  wire [28:0] _GEN_10; // @[Shift.scala 90:39]
  wire [28:0] _T_976; // @[Shift.scala 90:39]
  wire  _T_977; // @[Shift.scala 12:21]
  wire  _T_978; // @[Shift.scala 12:21]
  wire [1:0] _T_980; // @[Bitwise.scala 71:12]
  wire [30:0] _T_981; // @[Cat.scala 29:58]
  wire [30:0] _T_982; // @[Shift.scala 91:22]
  wire  _T_983; // @[Shift.scala 92:77]
  wire [29:0] _T_984; // @[Shift.scala 90:30]
  wire  _T_985; // @[Shift.scala 90:48]
  wire [29:0] _GEN_11; // @[Shift.scala 90:39]
  wire [29:0] _T_987; // @[Shift.scala 90:39]
  wire  _T_989; // @[Shift.scala 12:21]
  wire [30:0] _T_990; // @[Cat.scala 29:58]
  wire [30:0] _T_991; // @[Shift.scala 91:22]
  wire [30:0] _T_994; // @[Bitwise.scala 71:12]
  wire [30:0] _T_995; // @[Shift.scala 39:10]
  wire  _T_996; // @[convert.scala 55:31]
  wire  _T_997; // @[convert.scala 56:31]
  wire  _T_998; // @[convert.scala 57:31]
  wire  _T_999; // @[convert.scala 58:31]
  wire [27:0] _T_1000; // @[convert.scala 59:69]
  wire  _T_1001; // @[convert.scala 59:81]
  wire  _T_1002; // @[convert.scala 59:50]
  wire  _T_1004; // @[convert.scala 60:81]
  wire  _T_1005; // @[convert.scala 61:44]
  wire  _T_1006; // @[convert.scala 61:52]
  wire  _T_1007; // @[convert.scala 61:36]
  wire  _T_1008; // @[convert.scala 62:63]
  wire  _T_1009; // @[convert.scala 62:103]
  wire  _T_1010; // @[convert.scala 62:60]
  wire [27:0] _GEN_12; // @[convert.scala 63:56]
  wire [27:0] _T_1013; // @[convert.scala 63:56]
  wire [28:0] _T_1014; // @[Cat.scala 29:58]
  wire [28:0] _T_1016; // @[Mux.scala 87:16]
  assign _T_1 = io_A[28]; // @[convert.scala 18:24]
  assign _T_2 = io_A[27]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[27:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[26:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[26:11]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[15:8]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[7:4]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9[3:2]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10 != 2'h0; // @[LZD.scala 39:14]
  assign _T_12 = _T_10[1]; // @[LZD.scala 39:21]
  assign _T_13 = _T_10[0]; // @[LZD.scala 39:30]
  assign _T_14 = ~ _T_13; // @[LZD.scala 39:27]
  assign _T_15 = _T_12 | _T_14; // @[LZD.scala 39:25]
  assign _T_16 = {_T_11,_T_15}; // @[Cat.scala 29:58]
  assign _T_17 = _T_9[1:0]; // @[LZD.scala 44:32]
  assign _T_18 = _T_17 != 2'h0; // @[LZD.scala 39:14]
  assign _T_19 = _T_17[1]; // @[LZD.scala 39:21]
  assign _T_20 = _T_17[0]; // @[LZD.scala 39:30]
  assign _T_21 = ~ _T_20; // @[LZD.scala 39:27]
  assign _T_22 = _T_19 | _T_21; // @[LZD.scala 39:25]
  assign _T_23 = {_T_18,_T_22}; // @[Cat.scala 29:58]
  assign _T_24 = _T_16[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23[1]; // @[Shift.scala 12:21]
  assign _T_26 = _T_24 | _T_25; // @[LZD.scala 49:16]
  assign _T_27 = ~ _T_25; // @[LZD.scala 49:27]
  assign _T_28 = _T_24 | _T_27; // @[LZD.scala 49:25]
  assign _T_29 = _T_16[0:0]; // @[LZD.scala 49:47]
  assign _T_30 = _T_23[0:0]; // @[LZD.scala 49:59]
  assign _T_31 = _T_24 ? _T_29 : _T_30; // @[LZD.scala 49:35]
  assign _T_33 = {_T_26,_T_28,_T_31}; // @[Cat.scala 29:58]
  assign _T_34 = _T_8[3:0]; // @[LZD.scala 44:32]
  assign _T_35 = _T_34[3:2]; // @[LZD.scala 43:32]
  assign _T_36 = _T_35 != 2'h0; // @[LZD.scala 39:14]
  assign _T_37 = _T_35[1]; // @[LZD.scala 39:21]
  assign _T_38 = _T_35[0]; // @[LZD.scala 39:30]
  assign _T_39 = ~ _T_38; // @[LZD.scala 39:27]
  assign _T_40 = _T_37 | _T_39; // @[LZD.scala 39:25]
  assign _T_41 = {_T_36,_T_40}; // @[Cat.scala 29:58]
  assign _T_42 = _T_34[1:0]; // @[LZD.scala 44:32]
  assign _T_43 = _T_42 != 2'h0; // @[LZD.scala 39:14]
  assign _T_44 = _T_42[1]; // @[LZD.scala 39:21]
  assign _T_45 = _T_42[0]; // @[LZD.scala 39:30]
  assign _T_46 = ~ _T_45; // @[LZD.scala 39:27]
  assign _T_47 = _T_44 | _T_46; // @[LZD.scala 39:25]
  assign _T_48 = {_T_43,_T_47}; // @[Cat.scala 29:58]
  assign _T_49 = _T_41[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48[1]; // @[Shift.scala 12:21]
  assign _T_51 = _T_49 | _T_50; // @[LZD.scala 49:16]
  assign _T_52 = ~ _T_50; // @[LZD.scala 49:27]
  assign _T_53 = _T_49 | _T_52; // @[LZD.scala 49:25]
  assign _T_54 = _T_41[0:0]; // @[LZD.scala 49:47]
  assign _T_55 = _T_48[0:0]; // @[LZD.scala 49:59]
  assign _T_56 = _T_49 ? _T_54 : _T_55; // @[LZD.scala 49:35]
  assign _T_58 = {_T_51,_T_53,_T_56}; // @[Cat.scala 29:58]
  assign _T_59 = _T_33[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58[2]; // @[Shift.scala 12:21]
  assign _T_61 = _T_59 | _T_60; // @[LZD.scala 49:16]
  assign _T_62 = ~ _T_60; // @[LZD.scala 49:27]
  assign _T_63 = _T_59 | _T_62; // @[LZD.scala 49:25]
  assign _T_64 = _T_33[1:0]; // @[LZD.scala 49:47]
  assign _T_65 = _T_58[1:0]; // @[LZD.scala 49:59]
  assign _T_66 = _T_59 ? _T_64 : _T_65; // @[LZD.scala 49:35]
  assign _T_68 = {_T_61,_T_63,_T_66}; // @[Cat.scala 29:58]
  assign _T_69 = _T_7[7:0]; // @[LZD.scala 44:32]
  assign _T_70 = _T_69[7:4]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70[3:2]; // @[LZD.scala 43:32]
  assign _T_72 = _T_71 != 2'h0; // @[LZD.scala 39:14]
  assign _T_73 = _T_71[1]; // @[LZD.scala 39:21]
  assign _T_74 = _T_71[0]; // @[LZD.scala 39:30]
  assign _T_75 = ~ _T_74; // @[LZD.scala 39:27]
  assign _T_76 = _T_73 | _T_75; // @[LZD.scala 39:25]
  assign _T_77 = {_T_72,_T_76}; // @[Cat.scala 29:58]
  assign _T_78 = _T_70[1:0]; // @[LZD.scala 44:32]
  assign _T_79 = _T_78 != 2'h0; // @[LZD.scala 39:14]
  assign _T_80 = _T_78[1]; // @[LZD.scala 39:21]
  assign _T_81 = _T_78[0]; // @[LZD.scala 39:30]
  assign _T_82 = ~ _T_81; // @[LZD.scala 39:27]
  assign _T_83 = _T_80 | _T_82; // @[LZD.scala 39:25]
  assign _T_84 = {_T_79,_T_83}; // @[Cat.scala 29:58]
  assign _T_85 = _T_77[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84[1]; // @[Shift.scala 12:21]
  assign _T_87 = _T_85 | _T_86; // @[LZD.scala 49:16]
  assign _T_88 = ~ _T_86; // @[LZD.scala 49:27]
  assign _T_89 = _T_85 | _T_88; // @[LZD.scala 49:25]
  assign _T_90 = _T_77[0:0]; // @[LZD.scala 49:47]
  assign _T_91 = _T_84[0:0]; // @[LZD.scala 49:59]
  assign _T_92 = _T_85 ? _T_90 : _T_91; // @[LZD.scala 49:35]
  assign _T_94 = {_T_87,_T_89,_T_92}; // @[Cat.scala 29:58]
  assign _T_95 = _T_69[3:0]; // @[LZD.scala 44:32]
  assign _T_96 = _T_95[3:2]; // @[LZD.scala 43:32]
  assign _T_97 = _T_96 != 2'h0; // @[LZD.scala 39:14]
  assign _T_98 = _T_96[1]; // @[LZD.scala 39:21]
  assign _T_99 = _T_96[0]; // @[LZD.scala 39:30]
  assign _T_100 = ~ _T_99; // @[LZD.scala 39:27]
  assign _T_101 = _T_98 | _T_100; // @[LZD.scala 39:25]
  assign _T_102 = {_T_97,_T_101}; // @[Cat.scala 29:58]
  assign _T_103 = _T_95[1:0]; // @[LZD.scala 44:32]
  assign _T_104 = _T_103 != 2'h0; // @[LZD.scala 39:14]
  assign _T_105 = _T_103[1]; // @[LZD.scala 39:21]
  assign _T_106 = _T_103[0]; // @[LZD.scala 39:30]
  assign _T_107 = ~ _T_106; // @[LZD.scala 39:27]
  assign _T_108 = _T_105 | _T_107; // @[LZD.scala 39:25]
  assign _T_109 = {_T_104,_T_108}; // @[Cat.scala 29:58]
  assign _T_110 = _T_102[1]; // @[Shift.scala 12:21]
  assign _T_111 = _T_109[1]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110 | _T_111; // @[LZD.scala 49:16]
  assign _T_113 = ~ _T_111; // @[LZD.scala 49:27]
  assign _T_114 = _T_110 | _T_113; // @[LZD.scala 49:25]
  assign _T_115 = _T_102[0:0]; // @[LZD.scala 49:47]
  assign _T_116 = _T_109[0:0]; // @[LZD.scala 49:59]
  assign _T_117 = _T_110 ? _T_115 : _T_116; // @[LZD.scala 49:35]
  assign _T_119 = {_T_112,_T_114,_T_117}; // @[Cat.scala 29:58]
  assign _T_120 = _T_94[2]; // @[Shift.scala 12:21]
  assign _T_121 = _T_119[2]; // @[Shift.scala 12:21]
  assign _T_122 = _T_120 | _T_121; // @[LZD.scala 49:16]
  assign _T_123 = ~ _T_121; // @[LZD.scala 49:27]
  assign _T_124 = _T_120 | _T_123; // @[LZD.scala 49:25]
  assign _T_125 = _T_94[1:0]; // @[LZD.scala 49:47]
  assign _T_126 = _T_119[1:0]; // @[LZD.scala 49:59]
  assign _T_127 = _T_120 ? _T_125 : _T_126; // @[LZD.scala 49:35]
  assign _T_129 = {_T_122,_T_124,_T_127}; // @[Cat.scala 29:58]
  assign _T_130 = _T_68[3]; // @[Shift.scala 12:21]
  assign _T_131 = _T_129[3]; // @[Shift.scala 12:21]
  assign _T_132 = _T_130 | _T_131; // @[LZD.scala 49:16]
  assign _T_133 = ~ _T_131; // @[LZD.scala 49:27]
  assign _T_134 = _T_130 | _T_133; // @[LZD.scala 49:25]
  assign _T_135 = _T_68[2:0]; // @[LZD.scala 49:47]
  assign _T_136 = _T_129[2:0]; // @[LZD.scala 49:59]
  assign _T_137 = _T_130 ? _T_135 : _T_136; // @[LZD.scala 49:35]
  assign _T_139 = {_T_132,_T_134,_T_137}; // @[Cat.scala 29:58]
  assign _T_140 = _T_6[10:0]; // @[LZD.scala 44:32]
  assign _T_141 = _T_140[10:3]; // @[LZD.scala 43:32]
  assign _T_142 = _T_141[7:4]; // @[LZD.scala 43:32]
  assign _T_143 = _T_142[3:2]; // @[LZD.scala 43:32]
  assign _T_144 = _T_143 != 2'h0; // @[LZD.scala 39:14]
  assign _T_145 = _T_143[1]; // @[LZD.scala 39:21]
  assign _T_146 = _T_143[0]; // @[LZD.scala 39:30]
  assign _T_147 = ~ _T_146; // @[LZD.scala 39:27]
  assign _T_148 = _T_145 | _T_147; // @[LZD.scala 39:25]
  assign _T_149 = {_T_144,_T_148}; // @[Cat.scala 29:58]
  assign _T_150 = _T_142[1:0]; // @[LZD.scala 44:32]
  assign _T_151 = _T_150 != 2'h0; // @[LZD.scala 39:14]
  assign _T_152 = _T_150[1]; // @[LZD.scala 39:21]
  assign _T_153 = _T_150[0]; // @[LZD.scala 39:30]
  assign _T_154 = ~ _T_153; // @[LZD.scala 39:27]
  assign _T_155 = _T_152 | _T_154; // @[LZD.scala 39:25]
  assign _T_156 = {_T_151,_T_155}; // @[Cat.scala 29:58]
  assign _T_157 = _T_149[1]; // @[Shift.scala 12:21]
  assign _T_158 = _T_156[1]; // @[Shift.scala 12:21]
  assign _T_159 = _T_157 | _T_158; // @[LZD.scala 49:16]
  assign _T_160 = ~ _T_158; // @[LZD.scala 49:27]
  assign _T_161 = _T_157 | _T_160; // @[LZD.scala 49:25]
  assign _T_162 = _T_149[0:0]; // @[LZD.scala 49:47]
  assign _T_163 = _T_156[0:0]; // @[LZD.scala 49:59]
  assign _T_164 = _T_157 ? _T_162 : _T_163; // @[LZD.scala 49:35]
  assign _T_166 = {_T_159,_T_161,_T_164}; // @[Cat.scala 29:58]
  assign _T_167 = _T_141[3:0]; // @[LZD.scala 44:32]
  assign _T_168 = _T_167[3:2]; // @[LZD.scala 43:32]
  assign _T_169 = _T_168 != 2'h0; // @[LZD.scala 39:14]
  assign _T_170 = _T_168[1]; // @[LZD.scala 39:21]
  assign _T_171 = _T_168[0]; // @[LZD.scala 39:30]
  assign _T_172 = ~ _T_171; // @[LZD.scala 39:27]
  assign _T_173 = _T_170 | _T_172; // @[LZD.scala 39:25]
  assign _T_174 = {_T_169,_T_173}; // @[Cat.scala 29:58]
  assign _T_175 = _T_167[1:0]; // @[LZD.scala 44:32]
  assign _T_176 = _T_175 != 2'h0; // @[LZD.scala 39:14]
  assign _T_177 = _T_175[1]; // @[LZD.scala 39:21]
  assign _T_178 = _T_175[0]; // @[LZD.scala 39:30]
  assign _T_179 = ~ _T_178; // @[LZD.scala 39:27]
  assign _T_180 = _T_177 | _T_179; // @[LZD.scala 39:25]
  assign _T_181 = {_T_176,_T_180}; // @[Cat.scala 29:58]
  assign _T_182 = _T_174[1]; // @[Shift.scala 12:21]
  assign _T_183 = _T_181[1]; // @[Shift.scala 12:21]
  assign _T_184 = _T_182 | _T_183; // @[LZD.scala 49:16]
  assign _T_185 = ~ _T_183; // @[LZD.scala 49:27]
  assign _T_186 = _T_182 | _T_185; // @[LZD.scala 49:25]
  assign _T_187 = _T_174[0:0]; // @[LZD.scala 49:47]
  assign _T_188 = _T_181[0:0]; // @[LZD.scala 49:59]
  assign _T_189 = _T_182 ? _T_187 : _T_188; // @[LZD.scala 49:35]
  assign _T_191 = {_T_184,_T_186,_T_189}; // @[Cat.scala 29:58]
  assign _T_192 = _T_166[2]; // @[Shift.scala 12:21]
  assign _T_193 = _T_191[2]; // @[Shift.scala 12:21]
  assign _T_194 = _T_192 | _T_193; // @[LZD.scala 49:16]
  assign _T_195 = ~ _T_193; // @[LZD.scala 49:27]
  assign _T_196 = _T_192 | _T_195; // @[LZD.scala 49:25]
  assign _T_197 = _T_166[1:0]; // @[LZD.scala 49:47]
  assign _T_198 = _T_191[1:0]; // @[LZD.scala 49:59]
  assign _T_199 = _T_192 ? _T_197 : _T_198; // @[LZD.scala 49:35]
  assign _T_201 = {_T_194,_T_196,_T_199}; // @[Cat.scala 29:58]
  assign _T_202 = _T_140[2:0]; // @[LZD.scala 44:32]
  assign _T_203 = _T_202[2:1]; // @[LZD.scala 43:32]
  assign _T_204 = _T_203 != 2'h0; // @[LZD.scala 39:14]
  assign _T_205 = _T_203[1]; // @[LZD.scala 39:21]
  assign _T_206 = _T_203[0]; // @[LZD.scala 39:30]
  assign _T_207 = ~ _T_206; // @[LZD.scala 39:27]
  assign _T_208 = _T_205 | _T_207; // @[LZD.scala 39:25]
  assign _T_209 = {_T_204,_T_208}; // @[Cat.scala 29:58]
  assign _T_210 = _T_202[0:0]; // @[LZD.scala 44:32]
  assign _T_212 = _T_209[1]; // @[Shift.scala 12:21]
  assign _T_214 = _T_209[0:0]; // @[LZD.scala 55:32]
  assign _T_215 = _T_212 ? _T_214 : _T_210; // @[LZD.scala 55:20]
  assign _T_217 = _T_201[3]; // @[Shift.scala 12:21]
  assign _T_219 = {1'h1,_T_212,_T_215}; // @[Cat.scala 29:58]
  assign _T_220 = _T_201[2:0]; // @[LZD.scala 55:32]
  assign _T_221 = _T_217 ? _T_220 : _T_219; // @[LZD.scala 55:20]
  assign _T_222 = {_T_217,_T_221}; // @[Cat.scala 29:58]
  assign _T_223 = _T_139[4]; // @[Shift.scala 12:21]
  assign _T_225 = _T_139[3:0]; // @[LZD.scala 55:32]
  assign _T_226 = _T_223 ? _T_225 : _T_222; // @[LZD.scala 55:20]
  assign _T_227 = {_T_223,_T_226}; // @[Cat.scala 29:58]
  assign _T_228 = ~ _T_227; // @[convert.scala 21:22]
  assign _T_229 = io_A[25:0]; // @[convert.scala 22:36]
  assign _T_230 = _T_228 < 5'h1a; // @[Shift.scala 16:24]
  assign _T_232 = _T_228[4]; // @[Shift.scala 12:21]
  assign _T_233 = _T_229[9:0]; // @[Shift.scala 64:52]
  assign _T_235 = {_T_233,16'h0}; // @[Cat.scala 29:58]
  assign _T_236 = _T_232 ? _T_235 : _T_229; // @[Shift.scala 64:27]
  assign _T_237 = _T_228[3:0]; // @[Shift.scala 66:70]
  assign _T_238 = _T_237[3]; // @[Shift.scala 12:21]
  assign _T_239 = _T_236[17:0]; // @[Shift.scala 64:52]
  assign _T_241 = {_T_239,8'h0}; // @[Cat.scala 29:58]
  assign _T_242 = _T_238 ? _T_241 : _T_236; // @[Shift.scala 64:27]
  assign _T_243 = _T_237[2:0]; // @[Shift.scala 66:70]
  assign _T_244 = _T_243[2]; // @[Shift.scala 12:21]
  assign _T_245 = _T_242[21:0]; // @[Shift.scala 64:52]
  assign _T_247 = {_T_245,4'h0}; // @[Cat.scala 29:58]
  assign _T_248 = _T_244 ? _T_247 : _T_242; // @[Shift.scala 64:27]
  assign _T_249 = _T_243[1:0]; // @[Shift.scala 66:70]
  assign _T_250 = _T_249[1]; // @[Shift.scala 12:21]
  assign _T_251 = _T_248[23:0]; // @[Shift.scala 64:52]
  assign _T_253 = {_T_251,2'h0}; // @[Cat.scala 29:58]
  assign _T_254 = _T_250 ? _T_253 : _T_248; // @[Shift.scala 64:27]
  assign _T_255 = _T_249[0:0]; // @[Shift.scala 66:70]
  assign _T_257 = _T_254[24:0]; // @[Shift.scala 64:52]
  assign _T_258 = {_T_257,1'h0}; // @[Cat.scala 29:58]
  assign _T_259 = _T_255 ? _T_258 : _T_254; // @[Shift.scala 64:27]
  assign _T_260 = _T_230 ? _T_259 : 26'h0; // @[Shift.scala 16:10]
  assign _T_261 = _T_260[25:23]; // @[convert.scala 23:34]
  assign decA_fraction = _T_260[22:0]; // @[convert.scala 24:34]
  assign _T_263 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_265 = _T_3 ? _T_228 : _T_227; // @[convert.scala 25:42]
  assign _T_268 = ~ _T_261; // @[convert.scala 26:67]
  assign _T_269 = _T_1 ? _T_268 : _T_261; // @[convert.scala 26:51]
  assign _T_270 = {_T_263,_T_265,_T_269}; // @[Cat.scala 29:58]
  assign _T_272 = io_A[27:0]; // @[convert.scala 29:56]
  assign _T_273 = _T_272 != 28'h0; // @[convert.scala 29:60]
  assign _T_274 = ~ _T_273; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_274; // @[convert.scala 29:39]
  assign _T_277 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_277 & _T_274; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_270); // @[convert.scala 32:24]
  assign _T_286 = io_B[28]; // @[convert.scala 18:24]
  assign _T_287 = io_B[27]; // @[convert.scala 18:40]
  assign _T_288 = _T_286 ^ _T_287; // @[convert.scala 18:36]
  assign _T_289 = io_B[27:1]; // @[convert.scala 19:24]
  assign _T_290 = io_B[26:0]; // @[convert.scala 19:43]
  assign _T_291 = _T_289 ^ _T_290; // @[convert.scala 19:39]
  assign _T_292 = _T_291[26:11]; // @[LZD.scala 43:32]
  assign _T_293 = _T_292[15:8]; // @[LZD.scala 43:32]
  assign _T_294 = _T_293[7:4]; // @[LZD.scala 43:32]
  assign _T_295 = _T_294[3:2]; // @[LZD.scala 43:32]
  assign _T_296 = _T_295 != 2'h0; // @[LZD.scala 39:14]
  assign _T_297 = _T_295[1]; // @[LZD.scala 39:21]
  assign _T_298 = _T_295[0]; // @[LZD.scala 39:30]
  assign _T_299 = ~ _T_298; // @[LZD.scala 39:27]
  assign _T_300 = _T_297 | _T_299; // @[LZD.scala 39:25]
  assign _T_301 = {_T_296,_T_300}; // @[Cat.scala 29:58]
  assign _T_302 = _T_294[1:0]; // @[LZD.scala 44:32]
  assign _T_303 = _T_302 != 2'h0; // @[LZD.scala 39:14]
  assign _T_304 = _T_302[1]; // @[LZD.scala 39:21]
  assign _T_305 = _T_302[0]; // @[LZD.scala 39:30]
  assign _T_306 = ~ _T_305; // @[LZD.scala 39:27]
  assign _T_307 = _T_304 | _T_306; // @[LZD.scala 39:25]
  assign _T_308 = {_T_303,_T_307}; // @[Cat.scala 29:58]
  assign _T_309 = _T_301[1]; // @[Shift.scala 12:21]
  assign _T_310 = _T_308[1]; // @[Shift.scala 12:21]
  assign _T_311 = _T_309 | _T_310; // @[LZD.scala 49:16]
  assign _T_312 = ~ _T_310; // @[LZD.scala 49:27]
  assign _T_313 = _T_309 | _T_312; // @[LZD.scala 49:25]
  assign _T_314 = _T_301[0:0]; // @[LZD.scala 49:47]
  assign _T_315 = _T_308[0:0]; // @[LZD.scala 49:59]
  assign _T_316 = _T_309 ? _T_314 : _T_315; // @[LZD.scala 49:35]
  assign _T_318 = {_T_311,_T_313,_T_316}; // @[Cat.scala 29:58]
  assign _T_319 = _T_293[3:0]; // @[LZD.scala 44:32]
  assign _T_320 = _T_319[3:2]; // @[LZD.scala 43:32]
  assign _T_321 = _T_320 != 2'h0; // @[LZD.scala 39:14]
  assign _T_322 = _T_320[1]; // @[LZD.scala 39:21]
  assign _T_323 = _T_320[0]; // @[LZD.scala 39:30]
  assign _T_324 = ~ _T_323; // @[LZD.scala 39:27]
  assign _T_325 = _T_322 | _T_324; // @[LZD.scala 39:25]
  assign _T_326 = {_T_321,_T_325}; // @[Cat.scala 29:58]
  assign _T_327 = _T_319[1:0]; // @[LZD.scala 44:32]
  assign _T_328 = _T_327 != 2'h0; // @[LZD.scala 39:14]
  assign _T_329 = _T_327[1]; // @[LZD.scala 39:21]
  assign _T_330 = _T_327[0]; // @[LZD.scala 39:30]
  assign _T_331 = ~ _T_330; // @[LZD.scala 39:27]
  assign _T_332 = _T_329 | _T_331; // @[LZD.scala 39:25]
  assign _T_333 = {_T_328,_T_332}; // @[Cat.scala 29:58]
  assign _T_334 = _T_326[1]; // @[Shift.scala 12:21]
  assign _T_335 = _T_333[1]; // @[Shift.scala 12:21]
  assign _T_336 = _T_334 | _T_335; // @[LZD.scala 49:16]
  assign _T_337 = ~ _T_335; // @[LZD.scala 49:27]
  assign _T_338 = _T_334 | _T_337; // @[LZD.scala 49:25]
  assign _T_339 = _T_326[0:0]; // @[LZD.scala 49:47]
  assign _T_340 = _T_333[0:0]; // @[LZD.scala 49:59]
  assign _T_341 = _T_334 ? _T_339 : _T_340; // @[LZD.scala 49:35]
  assign _T_343 = {_T_336,_T_338,_T_341}; // @[Cat.scala 29:58]
  assign _T_344 = _T_318[2]; // @[Shift.scala 12:21]
  assign _T_345 = _T_343[2]; // @[Shift.scala 12:21]
  assign _T_346 = _T_344 | _T_345; // @[LZD.scala 49:16]
  assign _T_347 = ~ _T_345; // @[LZD.scala 49:27]
  assign _T_348 = _T_344 | _T_347; // @[LZD.scala 49:25]
  assign _T_349 = _T_318[1:0]; // @[LZD.scala 49:47]
  assign _T_350 = _T_343[1:0]; // @[LZD.scala 49:59]
  assign _T_351 = _T_344 ? _T_349 : _T_350; // @[LZD.scala 49:35]
  assign _T_353 = {_T_346,_T_348,_T_351}; // @[Cat.scala 29:58]
  assign _T_354 = _T_292[7:0]; // @[LZD.scala 44:32]
  assign _T_355 = _T_354[7:4]; // @[LZD.scala 43:32]
  assign _T_356 = _T_355[3:2]; // @[LZD.scala 43:32]
  assign _T_357 = _T_356 != 2'h0; // @[LZD.scala 39:14]
  assign _T_358 = _T_356[1]; // @[LZD.scala 39:21]
  assign _T_359 = _T_356[0]; // @[LZD.scala 39:30]
  assign _T_360 = ~ _T_359; // @[LZD.scala 39:27]
  assign _T_361 = _T_358 | _T_360; // @[LZD.scala 39:25]
  assign _T_362 = {_T_357,_T_361}; // @[Cat.scala 29:58]
  assign _T_363 = _T_355[1:0]; // @[LZD.scala 44:32]
  assign _T_364 = _T_363 != 2'h0; // @[LZD.scala 39:14]
  assign _T_365 = _T_363[1]; // @[LZD.scala 39:21]
  assign _T_366 = _T_363[0]; // @[LZD.scala 39:30]
  assign _T_367 = ~ _T_366; // @[LZD.scala 39:27]
  assign _T_368 = _T_365 | _T_367; // @[LZD.scala 39:25]
  assign _T_369 = {_T_364,_T_368}; // @[Cat.scala 29:58]
  assign _T_370 = _T_362[1]; // @[Shift.scala 12:21]
  assign _T_371 = _T_369[1]; // @[Shift.scala 12:21]
  assign _T_372 = _T_370 | _T_371; // @[LZD.scala 49:16]
  assign _T_373 = ~ _T_371; // @[LZD.scala 49:27]
  assign _T_374 = _T_370 | _T_373; // @[LZD.scala 49:25]
  assign _T_375 = _T_362[0:0]; // @[LZD.scala 49:47]
  assign _T_376 = _T_369[0:0]; // @[LZD.scala 49:59]
  assign _T_377 = _T_370 ? _T_375 : _T_376; // @[LZD.scala 49:35]
  assign _T_379 = {_T_372,_T_374,_T_377}; // @[Cat.scala 29:58]
  assign _T_380 = _T_354[3:0]; // @[LZD.scala 44:32]
  assign _T_381 = _T_380[3:2]; // @[LZD.scala 43:32]
  assign _T_382 = _T_381 != 2'h0; // @[LZD.scala 39:14]
  assign _T_383 = _T_381[1]; // @[LZD.scala 39:21]
  assign _T_384 = _T_381[0]; // @[LZD.scala 39:30]
  assign _T_385 = ~ _T_384; // @[LZD.scala 39:27]
  assign _T_386 = _T_383 | _T_385; // @[LZD.scala 39:25]
  assign _T_387 = {_T_382,_T_386}; // @[Cat.scala 29:58]
  assign _T_388 = _T_380[1:0]; // @[LZD.scala 44:32]
  assign _T_389 = _T_388 != 2'h0; // @[LZD.scala 39:14]
  assign _T_390 = _T_388[1]; // @[LZD.scala 39:21]
  assign _T_391 = _T_388[0]; // @[LZD.scala 39:30]
  assign _T_392 = ~ _T_391; // @[LZD.scala 39:27]
  assign _T_393 = _T_390 | _T_392; // @[LZD.scala 39:25]
  assign _T_394 = {_T_389,_T_393}; // @[Cat.scala 29:58]
  assign _T_395 = _T_387[1]; // @[Shift.scala 12:21]
  assign _T_396 = _T_394[1]; // @[Shift.scala 12:21]
  assign _T_397 = _T_395 | _T_396; // @[LZD.scala 49:16]
  assign _T_398 = ~ _T_396; // @[LZD.scala 49:27]
  assign _T_399 = _T_395 | _T_398; // @[LZD.scala 49:25]
  assign _T_400 = _T_387[0:0]; // @[LZD.scala 49:47]
  assign _T_401 = _T_394[0:0]; // @[LZD.scala 49:59]
  assign _T_402 = _T_395 ? _T_400 : _T_401; // @[LZD.scala 49:35]
  assign _T_404 = {_T_397,_T_399,_T_402}; // @[Cat.scala 29:58]
  assign _T_405 = _T_379[2]; // @[Shift.scala 12:21]
  assign _T_406 = _T_404[2]; // @[Shift.scala 12:21]
  assign _T_407 = _T_405 | _T_406; // @[LZD.scala 49:16]
  assign _T_408 = ~ _T_406; // @[LZD.scala 49:27]
  assign _T_409 = _T_405 | _T_408; // @[LZD.scala 49:25]
  assign _T_410 = _T_379[1:0]; // @[LZD.scala 49:47]
  assign _T_411 = _T_404[1:0]; // @[LZD.scala 49:59]
  assign _T_412 = _T_405 ? _T_410 : _T_411; // @[LZD.scala 49:35]
  assign _T_414 = {_T_407,_T_409,_T_412}; // @[Cat.scala 29:58]
  assign _T_415 = _T_353[3]; // @[Shift.scala 12:21]
  assign _T_416 = _T_414[3]; // @[Shift.scala 12:21]
  assign _T_417 = _T_415 | _T_416; // @[LZD.scala 49:16]
  assign _T_418 = ~ _T_416; // @[LZD.scala 49:27]
  assign _T_419 = _T_415 | _T_418; // @[LZD.scala 49:25]
  assign _T_420 = _T_353[2:0]; // @[LZD.scala 49:47]
  assign _T_421 = _T_414[2:0]; // @[LZD.scala 49:59]
  assign _T_422 = _T_415 ? _T_420 : _T_421; // @[LZD.scala 49:35]
  assign _T_424 = {_T_417,_T_419,_T_422}; // @[Cat.scala 29:58]
  assign _T_425 = _T_291[10:0]; // @[LZD.scala 44:32]
  assign _T_426 = _T_425[10:3]; // @[LZD.scala 43:32]
  assign _T_427 = _T_426[7:4]; // @[LZD.scala 43:32]
  assign _T_428 = _T_427[3:2]; // @[LZD.scala 43:32]
  assign _T_429 = _T_428 != 2'h0; // @[LZD.scala 39:14]
  assign _T_430 = _T_428[1]; // @[LZD.scala 39:21]
  assign _T_431 = _T_428[0]; // @[LZD.scala 39:30]
  assign _T_432 = ~ _T_431; // @[LZD.scala 39:27]
  assign _T_433 = _T_430 | _T_432; // @[LZD.scala 39:25]
  assign _T_434 = {_T_429,_T_433}; // @[Cat.scala 29:58]
  assign _T_435 = _T_427[1:0]; // @[LZD.scala 44:32]
  assign _T_436 = _T_435 != 2'h0; // @[LZD.scala 39:14]
  assign _T_437 = _T_435[1]; // @[LZD.scala 39:21]
  assign _T_438 = _T_435[0]; // @[LZD.scala 39:30]
  assign _T_439 = ~ _T_438; // @[LZD.scala 39:27]
  assign _T_440 = _T_437 | _T_439; // @[LZD.scala 39:25]
  assign _T_441 = {_T_436,_T_440}; // @[Cat.scala 29:58]
  assign _T_442 = _T_434[1]; // @[Shift.scala 12:21]
  assign _T_443 = _T_441[1]; // @[Shift.scala 12:21]
  assign _T_444 = _T_442 | _T_443; // @[LZD.scala 49:16]
  assign _T_445 = ~ _T_443; // @[LZD.scala 49:27]
  assign _T_446 = _T_442 | _T_445; // @[LZD.scala 49:25]
  assign _T_447 = _T_434[0:0]; // @[LZD.scala 49:47]
  assign _T_448 = _T_441[0:0]; // @[LZD.scala 49:59]
  assign _T_449 = _T_442 ? _T_447 : _T_448; // @[LZD.scala 49:35]
  assign _T_451 = {_T_444,_T_446,_T_449}; // @[Cat.scala 29:58]
  assign _T_452 = _T_426[3:0]; // @[LZD.scala 44:32]
  assign _T_453 = _T_452[3:2]; // @[LZD.scala 43:32]
  assign _T_454 = _T_453 != 2'h0; // @[LZD.scala 39:14]
  assign _T_455 = _T_453[1]; // @[LZD.scala 39:21]
  assign _T_456 = _T_453[0]; // @[LZD.scala 39:30]
  assign _T_457 = ~ _T_456; // @[LZD.scala 39:27]
  assign _T_458 = _T_455 | _T_457; // @[LZD.scala 39:25]
  assign _T_459 = {_T_454,_T_458}; // @[Cat.scala 29:58]
  assign _T_460 = _T_452[1:0]; // @[LZD.scala 44:32]
  assign _T_461 = _T_460 != 2'h0; // @[LZD.scala 39:14]
  assign _T_462 = _T_460[1]; // @[LZD.scala 39:21]
  assign _T_463 = _T_460[0]; // @[LZD.scala 39:30]
  assign _T_464 = ~ _T_463; // @[LZD.scala 39:27]
  assign _T_465 = _T_462 | _T_464; // @[LZD.scala 39:25]
  assign _T_466 = {_T_461,_T_465}; // @[Cat.scala 29:58]
  assign _T_467 = _T_459[1]; // @[Shift.scala 12:21]
  assign _T_468 = _T_466[1]; // @[Shift.scala 12:21]
  assign _T_469 = _T_467 | _T_468; // @[LZD.scala 49:16]
  assign _T_470 = ~ _T_468; // @[LZD.scala 49:27]
  assign _T_471 = _T_467 | _T_470; // @[LZD.scala 49:25]
  assign _T_472 = _T_459[0:0]; // @[LZD.scala 49:47]
  assign _T_473 = _T_466[0:0]; // @[LZD.scala 49:59]
  assign _T_474 = _T_467 ? _T_472 : _T_473; // @[LZD.scala 49:35]
  assign _T_476 = {_T_469,_T_471,_T_474}; // @[Cat.scala 29:58]
  assign _T_477 = _T_451[2]; // @[Shift.scala 12:21]
  assign _T_478 = _T_476[2]; // @[Shift.scala 12:21]
  assign _T_479 = _T_477 | _T_478; // @[LZD.scala 49:16]
  assign _T_480 = ~ _T_478; // @[LZD.scala 49:27]
  assign _T_481 = _T_477 | _T_480; // @[LZD.scala 49:25]
  assign _T_482 = _T_451[1:0]; // @[LZD.scala 49:47]
  assign _T_483 = _T_476[1:0]; // @[LZD.scala 49:59]
  assign _T_484 = _T_477 ? _T_482 : _T_483; // @[LZD.scala 49:35]
  assign _T_486 = {_T_479,_T_481,_T_484}; // @[Cat.scala 29:58]
  assign _T_487 = _T_425[2:0]; // @[LZD.scala 44:32]
  assign _T_488 = _T_487[2:1]; // @[LZD.scala 43:32]
  assign _T_489 = _T_488 != 2'h0; // @[LZD.scala 39:14]
  assign _T_490 = _T_488[1]; // @[LZD.scala 39:21]
  assign _T_491 = _T_488[0]; // @[LZD.scala 39:30]
  assign _T_492 = ~ _T_491; // @[LZD.scala 39:27]
  assign _T_493 = _T_490 | _T_492; // @[LZD.scala 39:25]
  assign _T_494 = {_T_489,_T_493}; // @[Cat.scala 29:58]
  assign _T_495 = _T_487[0:0]; // @[LZD.scala 44:32]
  assign _T_497 = _T_494[1]; // @[Shift.scala 12:21]
  assign _T_499 = _T_494[0:0]; // @[LZD.scala 55:32]
  assign _T_500 = _T_497 ? _T_499 : _T_495; // @[LZD.scala 55:20]
  assign _T_502 = _T_486[3]; // @[Shift.scala 12:21]
  assign _T_504 = {1'h1,_T_497,_T_500}; // @[Cat.scala 29:58]
  assign _T_505 = _T_486[2:0]; // @[LZD.scala 55:32]
  assign _T_506 = _T_502 ? _T_505 : _T_504; // @[LZD.scala 55:20]
  assign _T_507 = {_T_502,_T_506}; // @[Cat.scala 29:58]
  assign _T_508 = _T_424[4]; // @[Shift.scala 12:21]
  assign _T_510 = _T_424[3:0]; // @[LZD.scala 55:32]
  assign _T_511 = _T_508 ? _T_510 : _T_507; // @[LZD.scala 55:20]
  assign _T_512 = {_T_508,_T_511}; // @[Cat.scala 29:58]
  assign _T_513 = ~ _T_512; // @[convert.scala 21:22]
  assign _T_514 = io_B[25:0]; // @[convert.scala 22:36]
  assign _T_515 = _T_513 < 5'h1a; // @[Shift.scala 16:24]
  assign _T_517 = _T_513[4]; // @[Shift.scala 12:21]
  assign _T_518 = _T_514[9:0]; // @[Shift.scala 64:52]
  assign _T_520 = {_T_518,16'h0}; // @[Cat.scala 29:58]
  assign _T_521 = _T_517 ? _T_520 : _T_514; // @[Shift.scala 64:27]
  assign _T_522 = _T_513[3:0]; // @[Shift.scala 66:70]
  assign _T_523 = _T_522[3]; // @[Shift.scala 12:21]
  assign _T_524 = _T_521[17:0]; // @[Shift.scala 64:52]
  assign _T_526 = {_T_524,8'h0}; // @[Cat.scala 29:58]
  assign _T_527 = _T_523 ? _T_526 : _T_521; // @[Shift.scala 64:27]
  assign _T_528 = _T_522[2:0]; // @[Shift.scala 66:70]
  assign _T_529 = _T_528[2]; // @[Shift.scala 12:21]
  assign _T_530 = _T_527[21:0]; // @[Shift.scala 64:52]
  assign _T_532 = {_T_530,4'h0}; // @[Cat.scala 29:58]
  assign _T_533 = _T_529 ? _T_532 : _T_527; // @[Shift.scala 64:27]
  assign _T_534 = _T_528[1:0]; // @[Shift.scala 66:70]
  assign _T_535 = _T_534[1]; // @[Shift.scala 12:21]
  assign _T_536 = _T_533[23:0]; // @[Shift.scala 64:52]
  assign _T_538 = {_T_536,2'h0}; // @[Cat.scala 29:58]
  assign _T_539 = _T_535 ? _T_538 : _T_533; // @[Shift.scala 64:27]
  assign _T_540 = _T_534[0:0]; // @[Shift.scala 66:70]
  assign _T_542 = _T_539[24:0]; // @[Shift.scala 64:52]
  assign _T_543 = {_T_542,1'h0}; // @[Cat.scala 29:58]
  assign _T_544 = _T_540 ? _T_543 : _T_539; // @[Shift.scala 64:27]
  assign _T_545 = _T_515 ? _T_544 : 26'h0; // @[Shift.scala 16:10]
  assign _T_546 = _T_545[25:23]; // @[convert.scala 23:34]
  assign decB_fraction = _T_545[22:0]; // @[convert.scala 24:34]
  assign _T_548 = _T_288 == 1'h0; // @[convert.scala 25:26]
  assign _T_550 = _T_288 ? _T_513 : _T_512; // @[convert.scala 25:42]
  assign _T_553 = ~ _T_546; // @[convert.scala 26:67]
  assign _T_554 = _T_286 ? _T_553 : _T_546; // @[convert.scala 26:51]
  assign _T_555 = {_T_548,_T_550,_T_554}; // @[Cat.scala 29:58]
  assign _T_557 = io_B[27:0]; // @[convert.scala 29:56]
  assign _T_558 = _T_557 != 28'h0; // @[convert.scala 29:60]
  assign _T_559 = ~ _T_558; // @[convert.scala 29:41]
  assign decB_isNaR = _T_286 & _T_559; // @[convert.scala 29:39]
  assign _T_562 = _T_286 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_562 & _T_559; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_555); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[PositAdder.scala 24:32]
  assign greaterSign = aGTb ? _T_1 : _T_286; // @[PositAdder.scala 25:24]
  assign smallerSign = aGTb ? _T_286 : _T_1; // @[PositAdder.scala 26:24]
  assign greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[PositAdder.scala 27:24]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[PositAdder.scala 28:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[PositAdder.scala 29:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[PositAdder.scala 30:24]
  assign _T_571 = $signed(greaterExp) - $signed(smallerExp); // @[PositAdder.scala 31:32]
  assign scale_diff = $signed(_T_571); // @[PositAdder.scala 31:32]
  assign _T_572 = ~ greaterSign; // @[PositAdder.scala 32:38]
  assign greaterSig = {greaterSign,_T_572,greaterFrac}; // @[Cat.scala 29:58]
  assign _T_574 = ~ smallerSign; // @[PositAdder.scala 33:38]
  assign _T_577 = {smallerSign,_T_574,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_578 = $unsigned(scale_diff); // @[PositAdder.scala 34:68]
  assign _T_579 = _T_578 < 9'h1c; // @[Shift.scala 39:24]
  assign _T_580 = _T_578[4:0]; // @[Shift.scala 40:44]
  assign _T_581 = _T_577[27:16]; // @[Shift.scala 90:30]
  assign _T_582 = _T_577[15:0]; // @[Shift.scala 90:48]
  assign _T_583 = _T_582 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{11'd0}, _T_583}; // @[Shift.scala 90:39]
  assign _T_584 = _T_581 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_585 = _T_580[4]; // @[Shift.scala 12:21]
  assign _T_586 = _T_577[27]; // @[Shift.scala 12:21]
  assign _T_588 = _T_586 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_589 = {_T_588,_T_584}; // @[Cat.scala 29:58]
  assign _T_590 = _T_585 ? _T_589 : _T_577; // @[Shift.scala 91:22]
  assign _T_591 = _T_580[3:0]; // @[Shift.scala 92:77]
  assign _T_592 = _T_590[27:8]; // @[Shift.scala 90:30]
  assign _T_593 = _T_590[7:0]; // @[Shift.scala 90:48]
  assign _T_594 = _T_593 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{19'd0}, _T_594}; // @[Shift.scala 90:39]
  assign _T_595 = _T_592 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_596 = _T_591[3]; // @[Shift.scala 12:21]
  assign _T_597 = _T_590[27]; // @[Shift.scala 12:21]
  assign _T_599 = _T_597 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_600 = {_T_599,_T_595}; // @[Cat.scala 29:58]
  assign _T_601 = _T_596 ? _T_600 : _T_590; // @[Shift.scala 91:22]
  assign _T_602 = _T_591[2:0]; // @[Shift.scala 92:77]
  assign _T_603 = _T_601[27:4]; // @[Shift.scala 90:30]
  assign _T_604 = _T_601[3:0]; // @[Shift.scala 90:48]
  assign _T_605 = _T_604 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{23'd0}, _T_605}; // @[Shift.scala 90:39]
  assign _T_606 = _T_603 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_607 = _T_602[2]; // @[Shift.scala 12:21]
  assign _T_608 = _T_601[27]; // @[Shift.scala 12:21]
  assign _T_610 = _T_608 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_611 = {_T_610,_T_606}; // @[Cat.scala 29:58]
  assign _T_612 = _T_607 ? _T_611 : _T_601; // @[Shift.scala 91:22]
  assign _T_613 = _T_602[1:0]; // @[Shift.scala 92:77]
  assign _T_614 = _T_612[27:2]; // @[Shift.scala 90:30]
  assign _T_615 = _T_612[1:0]; // @[Shift.scala 90:48]
  assign _T_616 = _T_615 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_3 = {{25'd0}, _T_616}; // @[Shift.scala 90:39]
  assign _T_617 = _T_614 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_618 = _T_613[1]; // @[Shift.scala 12:21]
  assign _T_619 = _T_612[27]; // @[Shift.scala 12:21]
  assign _T_621 = _T_619 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_622 = {_T_621,_T_617}; // @[Cat.scala 29:58]
  assign _T_623 = _T_618 ? _T_622 : _T_612; // @[Shift.scala 91:22]
  assign _T_624 = _T_613[0:0]; // @[Shift.scala 92:77]
  assign _T_625 = _T_623[27:1]; // @[Shift.scala 90:30]
  assign _T_626 = _T_623[0:0]; // @[Shift.scala 90:48]
  assign _GEN_4 = {{26'd0}, _T_626}; // @[Shift.scala 90:39]
  assign _T_628 = _T_625 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_630 = _T_623[27]; // @[Shift.scala 12:21]
  assign _T_631 = {_T_630,_T_628}; // @[Cat.scala 29:58]
  assign _T_632 = _T_624 ? _T_631 : _T_623; // @[Shift.scala 91:22]
  assign _T_635 = _T_586 ? 28'hfffffff : 28'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_579 ? _T_632 : _T_635; // @[Shift.scala 39:10]
  assign _T_636 = smallerSig[27:3]; // @[PositAdder.scala 35:45]
  assign rawSumSig = greaterSig + _T_636; // @[PositAdder.scala 35:32]
  assign _T_637 = _T_1 ^ _T_286; // @[PositAdder.scala 36:31]
  assign _T_638 = rawSumSig[25:25]; // @[PositAdder.scala 36:59]
  assign sumSign = _T_637 ^ _T_638; // @[PositAdder.scala 36:43]
  assign _T_639 = greaterSig + _T_636; // @[PositAdder.scala 37:48]
  assign _T_640 = smallerSig[2:0]; // @[PositAdder.scala 37:63]
  assign signSumSig = {sumSign,_T_639,_T_640}; // @[Cat.scala 29:58]
  assign _T_642 = signSumSig[28:1]; // @[PositAdder.scala 39:31]
  assign _T_643 = signSumSig[27:0]; // @[PositAdder.scala 39:66]
  assign sumXor = _T_642 ^ _T_643; // @[PositAdder.scala 39:49]
  assign _T_644 = sumXor[27:12]; // @[LZD.scala 43:32]
  assign _T_645 = _T_644[15:8]; // @[LZD.scala 43:32]
  assign _T_646 = _T_645[7:4]; // @[LZD.scala 43:32]
  assign _T_647 = _T_646[3:2]; // @[LZD.scala 43:32]
  assign _T_648 = _T_647 != 2'h0; // @[LZD.scala 39:14]
  assign _T_649 = _T_647[1]; // @[LZD.scala 39:21]
  assign _T_650 = _T_647[0]; // @[LZD.scala 39:30]
  assign _T_651 = ~ _T_650; // @[LZD.scala 39:27]
  assign _T_652 = _T_649 | _T_651; // @[LZD.scala 39:25]
  assign _T_653 = {_T_648,_T_652}; // @[Cat.scala 29:58]
  assign _T_654 = _T_646[1:0]; // @[LZD.scala 44:32]
  assign _T_655 = _T_654 != 2'h0; // @[LZD.scala 39:14]
  assign _T_656 = _T_654[1]; // @[LZD.scala 39:21]
  assign _T_657 = _T_654[0]; // @[LZD.scala 39:30]
  assign _T_658 = ~ _T_657; // @[LZD.scala 39:27]
  assign _T_659 = _T_656 | _T_658; // @[LZD.scala 39:25]
  assign _T_660 = {_T_655,_T_659}; // @[Cat.scala 29:58]
  assign _T_661 = _T_653[1]; // @[Shift.scala 12:21]
  assign _T_662 = _T_660[1]; // @[Shift.scala 12:21]
  assign _T_663 = _T_661 | _T_662; // @[LZD.scala 49:16]
  assign _T_664 = ~ _T_662; // @[LZD.scala 49:27]
  assign _T_665 = _T_661 | _T_664; // @[LZD.scala 49:25]
  assign _T_666 = _T_653[0:0]; // @[LZD.scala 49:47]
  assign _T_667 = _T_660[0:0]; // @[LZD.scala 49:59]
  assign _T_668 = _T_661 ? _T_666 : _T_667; // @[LZD.scala 49:35]
  assign _T_670 = {_T_663,_T_665,_T_668}; // @[Cat.scala 29:58]
  assign _T_671 = _T_645[3:0]; // @[LZD.scala 44:32]
  assign _T_672 = _T_671[3:2]; // @[LZD.scala 43:32]
  assign _T_673 = _T_672 != 2'h0; // @[LZD.scala 39:14]
  assign _T_674 = _T_672[1]; // @[LZD.scala 39:21]
  assign _T_675 = _T_672[0]; // @[LZD.scala 39:30]
  assign _T_676 = ~ _T_675; // @[LZD.scala 39:27]
  assign _T_677 = _T_674 | _T_676; // @[LZD.scala 39:25]
  assign _T_678 = {_T_673,_T_677}; // @[Cat.scala 29:58]
  assign _T_679 = _T_671[1:0]; // @[LZD.scala 44:32]
  assign _T_680 = _T_679 != 2'h0; // @[LZD.scala 39:14]
  assign _T_681 = _T_679[1]; // @[LZD.scala 39:21]
  assign _T_682 = _T_679[0]; // @[LZD.scala 39:30]
  assign _T_683 = ~ _T_682; // @[LZD.scala 39:27]
  assign _T_684 = _T_681 | _T_683; // @[LZD.scala 39:25]
  assign _T_685 = {_T_680,_T_684}; // @[Cat.scala 29:58]
  assign _T_686 = _T_678[1]; // @[Shift.scala 12:21]
  assign _T_687 = _T_685[1]; // @[Shift.scala 12:21]
  assign _T_688 = _T_686 | _T_687; // @[LZD.scala 49:16]
  assign _T_689 = ~ _T_687; // @[LZD.scala 49:27]
  assign _T_690 = _T_686 | _T_689; // @[LZD.scala 49:25]
  assign _T_691 = _T_678[0:0]; // @[LZD.scala 49:47]
  assign _T_692 = _T_685[0:0]; // @[LZD.scala 49:59]
  assign _T_693 = _T_686 ? _T_691 : _T_692; // @[LZD.scala 49:35]
  assign _T_695 = {_T_688,_T_690,_T_693}; // @[Cat.scala 29:58]
  assign _T_696 = _T_670[2]; // @[Shift.scala 12:21]
  assign _T_697 = _T_695[2]; // @[Shift.scala 12:21]
  assign _T_698 = _T_696 | _T_697; // @[LZD.scala 49:16]
  assign _T_699 = ~ _T_697; // @[LZD.scala 49:27]
  assign _T_700 = _T_696 | _T_699; // @[LZD.scala 49:25]
  assign _T_701 = _T_670[1:0]; // @[LZD.scala 49:47]
  assign _T_702 = _T_695[1:0]; // @[LZD.scala 49:59]
  assign _T_703 = _T_696 ? _T_701 : _T_702; // @[LZD.scala 49:35]
  assign _T_705 = {_T_698,_T_700,_T_703}; // @[Cat.scala 29:58]
  assign _T_706 = _T_644[7:0]; // @[LZD.scala 44:32]
  assign _T_707 = _T_706[7:4]; // @[LZD.scala 43:32]
  assign _T_708 = _T_707[3:2]; // @[LZD.scala 43:32]
  assign _T_709 = _T_708 != 2'h0; // @[LZD.scala 39:14]
  assign _T_710 = _T_708[1]; // @[LZD.scala 39:21]
  assign _T_711 = _T_708[0]; // @[LZD.scala 39:30]
  assign _T_712 = ~ _T_711; // @[LZD.scala 39:27]
  assign _T_713 = _T_710 | _T_712; // @[LZD.scala 39:25]
  assign _T_714 = {_T_709,_T_713}; // @[Cat.scala 29:58]
  assign _T_715 = _T_707[1:0]; // @[LZD.scala 44:32]
  assign _T_716 = _T_715 != 2'h0; // @[LZD.scala 39:14]
  assign _T_717 = _T_715[1]; // @[LZD.scala 39:21]
  assign _T_718 = _T_715[0]; // @[LZD.scala 39:30]
  assign _T_719 = ~ _T_718; // @[LZD.scala 39:27]
  assign _T_720 = _T_717 | _T_719; // @[LZD.scala 39:25]
  assign _T_721 = {_T_716,_T_720}; // @[Cat.scala 29:58]
  assign _T_722 = _T_714[1]; // @[Shift.scala 12:21]
  assign _T_723 = _T_721[1]; // @[Shift.scala 12:21]
  assign _T_724 = _T_722 | _T_723; // @[LZD.scala 49:16]
  assign _T_725 = ~ _T_723; // @[LZD.scala 49:27]
  assign _T_726 = _T_722 | _T_725; // @[LZD.scala 49:25]
  assign _T_727 = _T_714[0:0]; // @[LZD.scala 49:47]
  assign _T_728 = _T_721[0:0]; // @[LZD.scala 49:59]
  assign _T_729 = _T_722 ? _T_727 : _T_728; // @[LZD.scala 49:35]
  assign _T_731 = {_T_724,_T_726,_T_729}; // @[Cat.scala 29:58]
  assign _T_732 = _T_706[3:0]; // @[LZD.scala 44:32]
  assign _T_733 = _T_732[3:2]; // @[LZD.scala 43:32]
  assign _T_734 = _T_733 != 2'h0; // @[LZD.scala 39:14]
  assign _T_735 = _T_733[1]; // @[LZD.scala 39:21]
  assign _T_736 = _T_733[0]; // @[LZD.scala 39:30]
  assign _T_737 = ~ _T_736; // @[LZD.scala 39:27]
  assign _T_738 = _T_735 | _T_737; // @[LZD.scala 39:25]
  assign _T_739 = {_T_734,_T_738}; // @[Cat.scala 29:58]
  assign _T_740 = _T_732[1:0]; // @[LZD.scala 44:32]
  assign _T_741 = _T_740 != 2'h0; // @[LZD.scala 39:14]
  assign _T_742 = _T_740[1]; // @[LZD.scala 39:21]
  assign _T_743 = _T_740[0]; // @[LZD.scala 39:30]
  assign _T_744 = ~ _T_743; // @[LZD.scala 39:27]
  assign _T_745 = _T_742 | _T_744; // @[LZD.scala 39:25]
  assign _T_746 = {_T_741,_T_745}; // @[Cat.scala 29:58]
  assign _T_747 = _T_739[1]; // @[Shift.scala 12:21]
  assign _T_748 = _T_746[1]; // @[Shift.scala 12:21]
  assign _T_749 = _T_747 | _T_748; // @[LZD.scala 49:16]
  assign _T_750 = ~ _T_748; // @[LZD.scala 49:27]
  assign _T_751 = _T_747 | _T_750; // @[LZD.scala 49:25]
  assign _T_752 = _T_739[0:0]; // @[LZD.scala 49:47]
  assign _T_753 = _T_746[0:0]; // @[LZD.scala 49:59]
  assign _T_754 = _T_747 ? _T_752 : _T_753; // @[LZD.scala 49:35]
  assign _T_756 = {_T_749,_T_751,_T_754}; // @[Cat.scala 29:58]
  assign _T_757 = _T_731[2]; // @[Shift.scala 12:21]
  assign _T_758 = _T_756[2]; // @[Shift.scala 12:21]
  assign _T_759 = _T_757 | _T_758; // @[LZD.scala 49:16]
  assign _T_760 = ~ _T_758; // @[LZD.scala 49:27]
  assign _T_761 = _T_757 | _T_760; // @[LZD.scala 49:25]
  assign _T_762 = _T_731[1:0]; // @[LZD.scala 49:47]
  assign _T_763 = _T_756[1:0]; // @[LZD.scala 49:59]
  assign _T_764 = _T_757 ? _T_762 : _T_763; // @[LZD.scala 49:35]
  assign _T_766 = {_T_759,_T_761,_T_764}; // @[Cat.scala 29:58]
  assign _T_767 = _T_705[3]; // @[Shift.scala 12:21]
  assign _T_768 = _T_766[3]; // @[Shift.scala 12:21]
  assign _T_769 = _T_767 | _T_768; // @[LZD.scala 49:16]
  assign _T_770 = ~ _T_768; // @[LZD.scala 49:27]
  assign _T_771 = _T_767 | _T_770; // @[LZD.scala 49:25]
  assign _T_772 = _T_705[2:0]; // @[LZD.scala 49:47]
  assign _T_773 = _T_766[2:0]; // @[LZD.scala 49:59]
  assign _T_774 = _T_767 ? _T_772 : _T_773; // @[LZD.scala 49:35]
  assign _T_776 = {_T_769,_T_771,_T_774}; // @[Cat.scala 29:58]
  assign _T_777 = sumXor[11:0]; // @[LZD.scala 44:32]
  assign _T_778 = _T_777[11:4]; // @[LZD.scala 43:32]
  assign _T_779 = _T_778[7:4]; // @[LZD.scala 43:32]
  assign _T_780 = _T_779[3:2]; // @[LZD.scala 43:32]
  assign _T_781 = _T_780 != 2'h0; // @[LZD.scala 39:14]
  assign _T_782 = _T_780[1]; // @[LZD.scala 39:21]
  assign _T_783 = _T_780[0]; // @[LZD.scala 39:30]
  assign _T_784 = ~ _T_783; // @[LZD.scala 39:27]
  assign _T_785 = _T_782 | _T_784; // @[LZD.scala 39:25]
  assign _T_786 = {_T_781,_T_785}; // @[Cat.scala 29:58]
  assign _T_787 = _T_779[1:0]; // @[LZD.scala 44:32]
  assign _T_788 = _T_787 != 2'h0; // @[LZD.scala 39:14]
  assign _T_789 = _T_787[1]; // @[LZD.scala 39:21]
  assign _T_790 = _T_787[0]; // @[LZD.scala 39:30]
  assign _T_791 = ~ _T_790; // @[LZD.scala 39:27]
  assign _T_792 = _T_789 | _T_791; // @[LZD.scala 39:25]
  assign _T_793 = {_T_788,_T_792}; // @[Cat.scala 29:58]
  assign _T_794 = _T_786[1]; // @[Shift.scala 12:21]
  assign _T_795 = _T_793[1]; // @[Shift.scala 12:21]
  assign _T_796 = _T_794 | _T_795; // @[LZD.scala 49:16]
  assign _T_797 = ~ _T_795; // @[LZD.scala 49:27]
  assign _T_798 = _T_794 | _T_797; // @[LZD.scala 49:25]
  assign _T_799 = _T_786[0:0]; // @[LZD.scala 49:47]
  assign _T_800 = _T_793[0:0]; // @[LZD.scala 49:59]
  assign _T_801 = _T_794 ? _T_799 : _T_800; // @[LZD.scala 49:35]
  assign _T_803 = {_T_796,_T_798,_T_801}; // @[Cat.scala 29:58]
  assign _T_804 = _T_778[3:0]; // @[LZD.scala 44:32]
  assign _T_805 = _T_804[3:2]; // @[LZD.scala 43:32]
  assign _T_806 = _T_805 != 2'h0; // @[LZD.scala 39:14]
  assign _T_807 = _T_805[1]; // @[LZD.scala 39:21]
  assign _T_808 = _T_805[0]; // @[LZD.scala 39:30]
  assign _T_809 = ~ _T_808; // @[LZD.scala 39:27]
  assign _T_810 = _T_807 | _T_809; // @[LZD.scala 39:25]
  assign _T_811 = {_T_806,_T_810}; // @[Cat.scala 29:58]
  assign _T_812 = _T_804[1:0]; // @[LZD.scala 44:32]
  assign _T_813 = _T_812 != 2'h0; // @[LZD.scala 39:14]
  assign _T_814 = _T_812[1]; // @[LZD.scala 39:21]
  assign _T_815 = _T_812[0]; // @[LZD.scala 39:30]
  assign _T_816 = ~ _T_815; // @[LZD.scala 39:27]
  assign _T_817 = _T_814 | _T_816; // @[LZD.scala 39:25]
  assign _T_818 = {_T_813,_T_817}; // @[Cat.scala 29:58]
  assign _T_819 = _T_811[1]; // @[Shift.scala 12:21]
  assign _T_820 = _T_818[1]; // @[Shift.scala 12:21]
  assign _T_821 = _T_819 | _T_820; // @[LZD.scala 49:16]
  assign _T_822 = ~ _T_820; // @[LZD.scala 49:27]
  assign _T_823 = _T_819 | _T_822; // @[LZD.scala 49:25]
  assign _T_824 = _T_811[0:0]; // @[LZD.scala 49:47]
  assign _T_825 = _T_818[0:0]; // @[LZD.scala 49:59]
  assign _T_826 = _T_819 ? _T_824 : _T_825; // @[LZD.scala 49:35]
  assign _T_828 = {_T_821,_T_823,_T_826}; // @[Cat.scala 29:58]
  assign _T_829 = _T_803[2]; // @[Shift.scala 12:21]
  assign _T_830 = _T_828[2]; // @[Shift.scala 12:21]
  assign _T_831 = _T_829 | _T_830; // @[LZD.scala 49:16]
  assign _T_832 = ~ _T_830; // @[LZD.scala 49:27]
  assign _T_833 = _T_829 | _T_832; // @[LZD.scala 49:25]
  assign _T_834 = _T_803[1:0]; // @[LZD.scala 49:47]
  assign _T_835 = _T_828[1:0]; // @[LZD.scala 49:59]
  assign _T_836 = _T_829 ? _T_834 : _T_835; // @[LZD.scala 49:35]
  assign _T_838 = {_T_831,_T_833,_T_836}; // @[Cat.scala 29:58]
  assign _T_839 = _T_777[3:0]; // @[LZD.scala 44:32]
  assign _T_840 = _T_839[3:2]; // @[LZD.scala 43:32]
  assign _T_841 = _T_840 != 2'h0; // @[LZD.scala 39:14]
  assign _T_842 = _T_840[1]; // @[LZD.scala 39:21]
  assign _T_843 = _T_840[0]; // @[LZD.scala 39:30]
  assign _T_844 = ~ _T_843; // @[LZD.scala 39:27]
  assign _T_845 = _T_842 | _T_844; // @[LZD.scala 39:25]
  assign _T_846 = {_T_841,_T_845}; // @[Cat.scala 29:58]
  assign _T_847 = _T_839[1:0]; // @[LZD.scala 44:32]
  assign _T_848 = _T_847 != 2'h0; // @[LZD.scala 39:14]
  assign _T_849 = _T_847[1]; // @[LZD.scala 39:21]
  assign _T_850 = _T_847[0]; // @[LZD.scala 39:30]
  assign _T_851 = ~ _T_850; // @[LZD.scala 39:27]
  assign _T_852 = _T_849 | _T_851; // @[LZD.scala 39:25]
  assign _T_853 = {_T_848,_T_852}; // @[Cat.scala 29:58]
  assign _T_854 = _T_846[1]; // @[Shift.scala 12:21]
  assign _T_855 = _T_853[1]; // @[Shift.scala 12:21]
  assign _T_856 = _T_854 | _T_855; // @[LZD.scala 49:16]
  assign _T_857 = ~ _T_855; // @[LZD.scala 49:27]
  assign _T_858 = _T_854 | _T_857; // @[LZD.scala 49:25]
  assign _T_859 = _T_846[0:0]; // @[LZD.scala 49:47]
  assign _T_860 = _T_853[0:0]; // @[LZD.scala 49:59]
  assign _T_861 = _T_854 ? _T_859 : _T_860; // @[LZD.scala 49:35]
  assign _T_863 = {_T_856,_T_858,_T_861}; // @[Cat.scala 29:58]
  assign _T_864 = _T_838[3]; // @[Shift.scala 12:21]
  assign _T_866 = _T_838[2:0]; // @[LZD.scala 55:32]
  assign _T_867 = _T_864 ? _T_866 : _T_863; // @[LZD.scala 55:20]
  assign _T_868 = {_T_864,_T_867}; // @[Cat.scala 29:58]
  assign _T_869 = _T_776[4]; // @[Shift.scala 12:21]
  assign _T_871 = _T_776[3:0]; // @[LZD.scala 55:32]
  assign _T_872 = _T_869 ? _T_871 : _T_868; // @[LZD.scala 55:20]
  assign sumLZD = {_T_869,_T_872}; // @[Cat.scala 29:58]
  assign _T_873 = {1'h1,_T_869,_T_872}; // @[Cat.scala 29:58]
  assign _T_874 = $signed(_T_873); // @[PositAdder.scala 41:38]
  assign _T_876 = $signed(_T_874) + $signed(6'sh2); // @[PositAdder.scala 41:45]
  assign scaleBias = $signed(_T_876); // @[PositAdder.scala 41:45]
  assign _GEN_5 = {{3{scaleBias[5]}},scaleBias}; // @[PositAdder.scala 42:32]
  assign sumScale = $signed(greaterExp) + $signed(_GEN_5); // @[PositAdder.scala 42:32]
  assign overflow = $signed(sumScale) > $signed(10'shd8); // @[PositAdder.scala 43:30]
  assign normalShift = ~ sumLZD; // @[PositAdder.scala 44:22]
  assign _T_877 = signSumSig[26:0]; // @[PositAdder.scala 45:36]
  assign _T_878 = normalShift < 5'h1b; // @[Shift.scala 16:24]
  assign _T_880 = normalShift[4]; // @[Shift.scala 12:21]
  assign _T_881 = _T_877[10:0]; // @[Shift.scala 64:52]
  assign _T_883 = {_T_881,16'h0}; // @[Cat.scala 29:58]
  assign _T_884 = _T_880 ? _T_883 : _T_877; // @[Shift.scala 64:27]
  assign _T_885 = normalShift[3:0]; // @[Shift.scala 66:70]
  assign _T_886 = _T_885[3]; // @[Shift.scala 12:21]
  assign _T_887 = _T_884[18:0]; // @[Shift.scala 64:52]
  assign _T_889 = {_T_887,8'h0}; // @[Cat.scala 29:58]
  assign _T_890 = _T_886 ? _T_889 : _T_884; // @[Shift.scala 64:27]
  assign _T_891 = _T_885[2:0]; // @[Shift.scala 66:70]
  assign _T_892 = _T_891[2]; // @[Shift.scala 12:21]
  assign _T_893 = _T_890[22:0]; // @[Shift.scala 64:52]
  assign _T_895 = {_T_893,4'h0}; // @[Cat.scala 29:58]
  assign _T_896 = _T_892 ? _T_895 : _T_890; // @[Shift.scala 64:27]
  assign _T_897 = _T_891[1:0]; // @[Shift.scala 66:70]
  assign _T_898 = _T_897[1]; // @[Shift.scala 12:21]
  assign _T_899 = _T_896[24:0]; // @[Shift.scala 64:52]
  assign _T_901 = {_T_899,2'h0}; // @[Cat.scala 29:58]
  assign _T_902 = _T_898 ? _T_901 : _T_896; // @[Shift.scala 64:27]
  assign _T_903 = _T_897[0:0]; // @[Shift.scala 66:70]
  assign _T_905 = _T_902[25:0]; // @[Shift.scala 64:52]
  assign _T_906 = {_T_905,1'h0}; // @[Cat.scala 29:58]
  assign _T_907 = _T_903 ? _T_906 : _T_902; // @[Shift.scala 64:27]
  assign shiftSig = _T_878 ? _T_907 : 27'h0; // @[Shift.scala 16:10]
  assign _T_908 = overflow ? $signed(10'shd8) : $signed(sumScale); // @[PositAdder.scala 50:24]
  assign decS_fraction = shiftSig[26:4]; // @[PositAdder.scala 51:34]
  assign decS_isNaR = decA_isNaR | decB_isNaR; // @[PositAdder.scala 52:32]
  assign _T_911 = signSumSig != 29'h0; // @[PositAdder.scala 53:33]
  assign _T_912 = ~ _T_911; // @[PositAdder.scala 53:21]
  assign _T_913 = decA_isZero & decB_isZero; // @[PositAdder.scala 53:52]
  assign decS_isZero = _T_912 | _T_913; // @[PositAdder.scala 53:37]
  assign _T_915 = shiftSig[3:2]; // @[PositAdder.scala 54:33]
  assign _T_916 = shiftSig[1]; // @[PositAdder.scala 54:49]
  assign _T_917 = shiftSig[0]; // @[PositAdder.scala 54:63]
  assign _T_918 = _T_916 | _T_917; // @[PositAdder.scala 54:53]
  assign _GEN_6 = _T_908[8:0]; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  assign decS_scale = $signed(_GEN_6); // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  assign _T_921 = decS_scale[2:0]; // @[convert.scala 46:61]
  assign _T_922 = ~ _T_921; // @[convert.scala 46:52]
  assign _T_924 = sumSign ? _T_922 : _T_921; // @[convert.scala 46:42]
  assign _T_925 = decS_scale[8:3]; // @[convert.scala 48:34]
  assign _T_926 = _T_925[5:5]; // @[convert.scala 49:36]
  assign _T_928 = ~ _T_925; // @[convert.scala 50:36]
  assign _T_929 = $signed(_T_928); // @[convert.scala 50:36]
  assign _T_930 = _T_926 ? $signed(_T_929) : $signed(_T_925); // @[convert.scala 50:28]
  assign _T_931 = _T_926 ^ sumSign; // @[convert.scala 51:31]
  assign _T_932 = ~ _T_931; // @[convert.scala 52:43]
  assign _T_936 = {_T_932,_T_931,_T_924,decS_fraction,_T_915,_T_918}; // @[Cat.scala 29:58]
  assign _T_937 = $unsigned(_T_930); // @[Shift.scala 39:17]
  assign _T_938 = _T_937 < 6'h1f; // @[Shift.scala 39:24]
  assign _T_939 = _T_930[4:0]; // @[Shift.scala 40:44]
  assign _T_940 = _T_936[30:16]; // @[Shift.scala 90:30]
  assign _T_941 = _T_936[15:0]; // @[Shift.scala 90:48]
  assign _T_942 = _T_941 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{14'd0}, _T_942}; // @[Shift.scala 90:39]
  assign _T_943 = _T_940 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_944 = _T_939[4]; // @[Shift.scala 12:21]
  assign _T_945 = _T_936[30]; // @[Shift.scala 12:21]
  assign _T_947 = _T_945 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_948 = {_T_947,_T_943}; // @[Cat.scala 29:58]
  assign _T_949 = _T_944 ? _T_948 : _T_936; // @[Shift.scala 91:22]
  assign _T_950 = _T_939[3:0]; // @[Shift.scala 92:77]
  assign _T_951 = _T_949[30:8]; // @[Shift.scala 90:30]
  assign _T_952 = _T_949[7:0]; // @[Shift.scala 90:48]
  assign _T_953 = _T_952 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_8 = {{22'd0}, _T_953}; // @[Shift.scala 90:39]
  assign _T_954 = _T_951 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_955 = _T_950[3]; // @[Shift.scala 12:21]
  assign _T_956 = _T_949[30]; // @[Shift.scala 12:21]
  assign _T_958 = _T_956 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_959 = {_T_958,_T_954}; // @[Cat.scala 29:58]
  assign _T_960 = _T_955 ? _T_959 : _T_949; // @[Shift.scala 91:22]
  assign _T_961 = _T_950[2:0]; // @[Shift.scala 92:77]
  assign _T_962 = _T_960[30:4]; // @[Shift.scala 90:30]
  assign _T_963 = _T_960[3:0]; // @[Shift.scala 90:48]
  assign _T_964 = _T_963 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_9 = {{26'd0}, _T_964}; // @[Shift.scala 90:39]
  assign _T_965 = _T_962 | _GEN_9; // @[Shift.scala 90:39]
  assign _T_966 = _T_961[2]; // @[Shift.scala 12:21]
  assign _T_967 = _T_960[30]; // @[Shift.scala 12:21]
  assign _T_969 = _T_967 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_970 = {_T_969,_T_965}; // @[Cat.scala 29:58]
  assign _T_971 = _T_966 ? _T_970 : _T_960; // @[Shift.scala 91:22]
  assign _T_972 = _T_961[1:0]; // @[Shift.scala 92:77]
  assign _T_973 = _T_971[30:2]; // @[Shift.scala 90:30]
  assign _T_974 = _T_971[1:0]; // @[Shift.scala 90:48]
  assign _T_975 = _T_974 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_10 = {{28'd0}, _T_975}; // @[Shift.scala 90:39]
  assign _T_976 = _T_973 | _GEN_10; // @[Shift.scala 90:39]
  assign _T_977 = _T_972[1]; // @[Shift.scala 12:21]
  assign _T_978 = _T_971[30]; // @[Shift.scala 12:21]
  assign _T_980 = _T_978 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_981 = {_T_980,_T_976}; // @[Cat.scala 29:58]
  assign _T_982 = _T_977 ? _T_981 : _T_971; // @[Shift.scala 91:22]
  assign _T_983 = _T_972[0:0]; // @[Shift.scala 92:77]
  assign _T_984 = _T_982[30:1]; // @[Shift.scala 90:30]
  assign _T_985 = _T_982[0:0]; // @[Shift.scala 90:48]
  assign _GEN_11 = {{29'd0}, _T_985}; // @[Shift.scala 90:39]
  assign _T_987 = _T_984 | _GEN_11; // @[Shift.scala 90:39]
  assign _T_989 = _T_982[30]; // @[Shift.scala 12:21]
  assign _T_990 = {_T_989,_T_987}; // @[Cat.scala 29:58]
  assign _T_991 = _T_983 ? _T_990 : _T_982; // @[Shift.scala 91:22]
  assign _T_994 = _T_945 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 71:12]
  assign _T_995 = _T_938 ? _T_991 : _T_994; // @[Shift.scala 39:10]
  assign _T_996 = _T_995[3]; // @[convert.scala 55:31]
  assign _T_997 = _T_995[2]; // @[convert.scala 56:31]
  assign _T_998 = _T_995[1]; // @[convert.scala 57:31]
  assign _T_999 = _T_995[0]; // @[convert.scala 58:31]
  assign _T_1000 = _T_995[30:3]; // @[convert.scala 59:69]
  assign _T_1001 = _T_1000 != 28'h0; // @[convert.scala 59:81]
  assign _T_1002 = ~ _T_1001; // @[convert.scala 59:50]
  assign _T_1004 = _T_1000 == 28'hfffffff; // @[convert.scala 60:81]
  assign _T_1005 = _T_996 | _T_998; // @[convert.scala 61:44]
  assign _T_1006 = _T_1005 | _T_999; // @[convert.scala 61:52]
  assign _T_1007 = _T_997 & _T_1006; // @[convert.scala 61:36]
  assign _T_1008 = ~ _T_1004; // @[convert.scala 62:63]
  assign _T_1009 = _T_1008 & _T_1007; // @[convert.scala 62:103]
  assign _T_1010 = _T_1002 | _T_1009; // @[convert.scala 62:60]
  assign _GEN_12 = {{27'd0}, _T_1010}; // @[convert.scala 63:56]
  assign _T_1013 = _T_1000 + _GEN_12; // @[convert.scala 63:56]
  assign _T_1014 = {sumSign,_T_1013}; // @[Cat.scala 29:58]
  assign _T_1016 = decS_isZero ? 29'h0 : _T_1014; // @[Mux.scala 87:16]
  assign io_S = decS_isNaR ? 29'h10000000 : _T_1016; // @[PositAdder.scala 56:8]
endmodule
