module PositAdder13_1(
  input         clock,
  input         reset,
  input  [12:0] io_A,
  input  [12:0] io_B,
  output [12:0] io_S
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [10:0] _T_4; // @[convert.scala 19:24]
  wire [10:0] _T_5; // @[convert.scala 19:43]
  wire [10:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [2:0] _T_68; // @[LZD.scala 44:32]
  wire [1:0] _T_69; // @[LZD.scala 43:32]
  wire  _T_70; // @[LZD.scala 39:14]
  wire  _T_71; // @[LZD.scala 39:21]
  wire  _T_72; // @[LZD.scala 39:30]
  wire  _T_73; // @[LZD.scala 39:27]
  wire  _T_74; // @[LZD.scala 39:25]
  wire [1:0] _T_75; // @[Cat.scala 29:58]
  wire  _T_76; // @[LZD.scala 44:32]
  wire  _T_78; // @[Shift.scala 12:21]
  wire  _T_80; // @[LZD.scala 55:32]
  wire  _T_81; // @[LZD.scala 55:20]
  wire  _T_83; // @[Shift.scala 12:21]
  wire [2:0] _T_85; // @[Cat.scala 29:58]
  wire [2:0] _T_86; // @[LZD.scala 55:32]
  wire [2:0] _T_87; // @[LZD.scala 55:20]
  wire [3:0] _T_88; // @[Cat.scala 29:58]
  wire [3:0] _T_89; // @[convert.scala 21:22]
  wire [9:0] _T_90; // @[convert.scala 22:36]
  wire  _T_91; // @[Shift.scala 16:24]
  wire  _T_93; // @[Shift.scala 12:21]
  wire [1:0] _T_94; // @[Shift.scala 64:52]
  wire [9:0] _T_96; // @[Cat.scala 29:58]
  wire [9:0] _T_97; // @[Shift.scala 64:27]
  wire [2:0] _T_98; // @[Shift.scala 66:70]
  wire  _T_99; // @[Shift.scala 12:21]
  wire [5:0] _T_100; // @[Shift.scala 64:52]
  wire [9:0] _T_102; // @[Cat.scala 29:58]
  wire [9:0] _T_103; // @[Shift.scala 64:27]
  wire [1:0] _T_104; // @[Shift.scala 66:70]
  wire  _T_105; // @[Shift.scala 12:21]
  wire [7:0] _T_106; // @[Shift.scala 64:52]
  wire [9:0] _T_108; // @[Cat.scala 29:58]
  wire [9:0] _T_109; // @[Shift.scala 64:27]
  wire  _T_110; // @[Shift.scala 66:70]
  wire [8:0] _T_112; // @[Shift.scala 64:52]
  wire [9:0] _T_113; // @[Cat.scala 29:58]
  wire [9:0] _T_114; // @[Shift.scala 64:27]
  wire [9:0] _T_115; // @[Shift.scala 16:10]
  wire  _T_116; // @[convert.scala 23:34]
  wire [8:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_118; // @[convert.scala 25:26]
  wire [3:0] _T_120; // @[convert.scala 25:42]
  wire  _T_123; // @[convert.scala 26:67]
  wire  _T_124; // @[convert.scala 26:51]
  wire [5:0] _T_125; // @[Cat.scala 29:58]
  wire [11:0] _T_127; // @[convert.scala 29:56]
  wire  _T_128; // @[convert.scala 29:60]
  wire  _T_129; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_132; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_141; // @[convert.scala 18:24]
  wire  _T_142; // @[convert.scala 18:40]
  wire  _T_143; // @[convert.scala 18:36]
  wire [10:0] _T_144; // @[convert.scala 19:24]
  wire [10:0] _T_145; // @[convert.scala 19:43]
  wire [10:0] _T_146; // @[convert.scala 19:39]
  wire [7:0] _T_147; // @[LZD.scala 43:32]
  wire [3:0] _T_148; // @[LZD.scala 43:32]
  wire [1:0] _T_149; // @[LZD.scala 43:32]
  wire  _T_150; // @[LZD.scala 39:14]
  wire  _T_151; // @[LZD.scala 39:21]
  wire  _T_152; // @[LZD.scala 39:30]
  wire  _T_153; // @[LZD.scala 39:27]
  wire  _T_154; // @[LZD.scala 39:25]
  wire [1:0] _T_155; // @[Cat.scala 29:58]
  wire [1:0] _T_156; // @[LZD.scala 44:32]
  wire  _T_157; // @[LZD.scala 39:14]
  wire  _T_158; // @[LZD.scala 39:21]
  wire  _T_159; // @[LZD.scala 39:30]
  wire  _T_160; // @[LZD.scala 39:27]
  wire  _T_161; // @[LZD.scala 39:25]
  wire [1:0] _T_162; // @[Cat.scala 29:58]
  wire  _T_163; // @[Shift.scala 12:21]
  wire  _T_164; // @[Shift.scala 12:21]
  wire  _T_165; // @[LZD.scala 49:16]
  wire  _T_166; // @[LZD.scala 49:27]
  wire  _T_167; // @[LZD.scala 49:25]
  wire  _T_168; // @[LZD.scala 49:47]
  wire  _T_169; // @[LZD.scala 49:59]
  wire  _T_170; // @[LZD.scala 49:35]
  wire [2:0] _T_172; // @[Cat.scala 29:58]
  wire [3:0] _T_173; // @[LZD.scala 44:32]
  wire [1:0] _T_174; // @[LZD.scala 43:32]
  wire  _T_175; // @[LZD.scala 39:14]
  wire  _T_176; // @[LZD.scala 39:21]
  wire  _T_177; // @[LZD.scala 39:30]
  wire  _T_178; // @[LZD.scala 39:27]
  wire  _T_179; // @[LZD.scala 39:25]
  wire [1:0] _T_180; // @[Cat.scala 29:58]
  wire [1:0] _T_181; // @[LZD.scala 44:32]
  wire  _T_182; // @[LZD.scala 39:14]
  wire  _T_183; // @[LZD.scala 39:21]
  wire  _T_184; // @[LZD.scala 39:30]
  wire  _T_185; // @[LZD.scala 39:27]
  wire  _T_186; // @[LZD.scala 39:25]
  wire [1:0] _T_187; // @[Cat.scala 29:58]
  wire  _T_188; // @[Shift.scala 12:21]
  wire  _T_189; // @[Shift.scala 12:21]
  wire  _T_190; // @[LZD.scala 49:16]
  wire  _T_191; // @[LZD.scala 49:27]
  wire  _T_192; // @[LZD.scala 49:25]
  wire  _T_193; // @[LZD.scala 49:47]
  wire  _T_194; // @[LZD.scala 49:59]
  wire  _T_195; // @[LZD.scala 49:35]
  wire [2:0] _T_197; // @[Cat.scala 29:58]
  wire  _T_198; // @[Shift.scala 12:21]
  wire  _T_199; // @[Shift.scala 12:21]
  wire  _T_200; // @[LZD.scala 49:16]
  wire  _T_201; // @[LZD.scala 49:27]
  wire  _T_202; // @[LZD.scala 49:25]
  wire [1:0] _T_203; // @[LZD.scala 49:47]
  wire [1:0] _T_204; // @[LZD.scala 49:59]
  wire [1:0] _T_205; // @[LZD.scala 49:35]
  wire [3:0] _T_207; // @[Cat.scala 29:58]
  wire [2:0] _T_208; // @[LZD.scala 44:32]
  wire [1:0] _T_209; // @[LZD.scala 43:32]
  wire  _T_210; // @[LZD.scala 39:14]
  wire  _T_211; // @[LZD.scala 39:21]
  wire  _T_212; // @[LZD.scala 39:30]
  wire  _T_213; // @[LZD.scala 39:27]
  wire  _T_214; // @[LZD.scala 39:25]
  wire [1:0] _T_215; // @[Cat.scala 29:58]
  wire  _T_216; // @[LZD.scala 44:32]
  wire  _T_218; // @[Shift.scala 12:21]
  wire  _T_220; // @[LZD.scala 55:32]
  wire  _T_221; // @[LZD.scala 55:20]
  wire  _T_223; // @[Shift.scala 12:21]
  wire [2:0] _T_225; // @[Cat.scala 29:58]
  wire [2:0] _T_226; // @[LZD.scala 55:32]
  wire [2:0] _T_227; // @[LZD.scala 55:20]
  wire [3:0] _T_228; // @[Cat.scala 29:58]
  wire [3:0] _T_229; // @[convert.scala 21:22]
  wire [9:0] _T_230; // @[convert.scala 22:36]
  wire  _T_231; // @[Shift.scala 16:24]
  wire  _T_233; // @[Shift.scala 12:21]
  wire [1:0] _T_234; // @[Shift.scala 64:52]
  wire [9:0] _T_236; // @[Cat.scala 29:58]
  wire [9:0] _T_237; // @[Shift.scala 64:27]
  wire [2:0] _T_238; // @[Shift.scala 66:70]
  wire  _T_239; // @[Shift.scala 12:21]
  wire [5:0] _T_240; // @[Shift.scala 64:52]
  wire [9:0] _T_242; // @[Cat.scala 29:58]
  wire [9:0] _T_243; // @[Shift.scala 64:27]
  wire [1:0] _T_244; // @[Shift.scala 66:70]
  wire  _T_245; // @[Shift.scala 12:21]
  wire [7:0] _T_246; // @[Shift.scala 64:52]
  wire [9:0] _T_248; // @[Cat.scala 29:58]
  wire [9:0] _T_249; // @[Shift.scala 64:27]
  wire  _T_250; // @[Shift.scala 66:70]
  wire [8:0] _T_252; // @[Shift.scala 64:52]
  wire [9:0] _T_253; // @[Cat.scala 29:58]
  wire [9:0] _T_254; // @[Shift.scala 64:27]
  wire [9:0] _T_255; // @[Shift.scala 16:10]
  wire  _T_256; // @[convert.scala 23:34]
  wire [8:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_258; // @[convert.scala 25:26]
  wire [3:0] _T_260; // @[convert.scala 25:42]
  wire  _T_263; // @[convert.scala 26:67]
  wire  _T_264; // @[convert.scala 26:51]
  wire [5:0] _T_265; // @[Cat.scala 29:58]
  wire [11:0] _T_267; // @[convert.scala 29:56]
  wire  _T_268; // @[convert.scala 29:60]
  wire  _T_269; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_272; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[PositAdder.scala 24:32]
  wire  greaterSign; // @[PositAdder.scala 25:24]
  wire  smallerSign; // @[PositAdder.scala 26:24]
  wire [5:0] greaterExp; // @[PositAdder.scala 27:24]
  wire [5:0] smallerExp; // @[PositAdder.scala 28:24]
  wire [8:0] greaterFrac; // @[PositAdder.scala 29:24]
  wire [8:0] smallerFrac; // @[PositAdder.scala 30:24]
  wire [5:0] _T_281; // @[PositAdder.scala 31:32]
  wire [5:0] scale_diff; // @[PositAdder.scala 31:32]
  wire  _T_282; // @[PositAdder.scala 32:38]
  wire [10:0] greaterSig; // @[Cat.scala 29:58]
  wire  _T_284; // @[PositAdder.scala 33:38]
  wire [13:0] _T_287; // @[Cat.scala 29:58]
  wire [5:0] _T_288; // @[PositAdder.scala 34:68]
  wire  _T_289; // @[Shift.scala 39:24]
  wire [3:0] _T_290; // @[Shift.scala 40:44]
  wire [5:0] _T_291; // @[Shift.scala 90:30]
  wire [7:0] _T_292; // @[Shift.scala 90:48]
  wire  _T_293; // @[Shift.scala 90:57]
  wire [5:0] _GEN_0; // @[Shift.scala 90:39]
  wire [5:0] _T_294; // @[Shift.scala 90:39]
  wire  _T_295; // @[Shift.scala 12:21]
  wire  _T_296; // @[Shift.scala 12:21]
  wire [7:0] _T_298; // @[Bitwise.scala 71:12]
  wire [13:0] _T_299; // @[Cat.scala 29:58]
  wire [13:0] _T_300; // @[Shift.scala 91:22]
  wire [2:0] _T_301; // @[Shift.scala 92:77]
  wire [9:0] _T_302; // @[Shift.scala 90:30]
  wire [3:0] _T_303; // @[Shift.scala 90:48]
  wire  _T_304; // @[Shift.scala 90:57]
  wire [9:0] _GEN_1; // @[Shift.scala 90:39]
  wire [9:0] _T_305; // @[Shift.scala 90:39]
  wire  _T_306; // @[Shift.scala 12:21]
  wire  _T_307; // @[Shift.scala 12:21]
  wire [3:0] _T_309; // @[Bitwise.scala 71:12]
  wire [13:0] _T_310; // @[Cat.scala 29:58]
  wire [13:0] _T_311; // @[Shift.scala 91:22]
  wire [1:0] _T_312; // @[Shift.scala 92:77]
  wire [11:0] _T_313; // @[Shift.scala 90:30]
  wire [1:0] _T_314; // @[Shift.scala 90:48]
  wire  _T_315; // @[Shift.scala 90:57]
  wire [11:0] _GEN_2; // @[Shift.scala 90:39]
  wire [11:0] _T_316; // @[Shift.scala 90:39]
  wire  _T_317; // @[Shift.scala 12:21]
  wire  _T_318; // @[Shift.scala 12:21]
  wire [1:0] _T_320; // @[Bitwise.scala 71:12]
  wire [13:0] _T_321; // @[Cat.scala 29:58]
  wire [13:0] _T_322; // @[Shift.scala 91:22]
  wire  _T_323; // @[Shift.scala 92:77]
  wire [12:0] _T_324; // @[Shift.scala 90:30]
  wire  _T_325; // @[Shift.scala 90:48]
  wire [12:0] _GEN_3; // @[Shift.scala 90:39]
  wire [12:0] _T_327; // @[Shift.scala 90:39]
  wire  _T_329; // @[Shift.scala 12:21]
  wire [13:0] _T_330; // @[Cat.scala 29:58]
  wire [13:0] _T_331; // @[Shift.scala 91:22]
  wire [13:0] _T_334; // @[Bitwise.scala 71:12]
  wire [13:0] smallerSig; // @[Shift.scala 39:10]
  wire [10:0] _T_335; // @[PositAdder.scala 35:45]
  wire [11:0] rawSumSig; // @[PositAdder.scala 35:32]
  wire  _T_336; // @[PositAdder.scala 36:31]
  wire  _T_337; // @[PositAdder.scala 36:59]
  wire  sumSign; // @[PositAdder.scala 36:43]
  wire [10:0] _T_338; // @[PositAdder.scala 37:48]
  wire [2:0] _T_339; // @[PositAdder.scala 37:63]
  wire [14:0] signSumSig; // @[Cat.scala 29:58]
  wire [13:0] _T_341; // @[PositAdder.scala 39:31]
  wire [13:0] _T_342; // @[PositAdder.scala 39:66]
  wire [13:0] sumXor; // @[PositAdder.scala 39:49]
  wire [7:0] _T_343; // @[LZD.scala 43:32]
  wire [3:0] _T_344; // @[LZD.scala 43:32]
  wire [1:0] _T_345; // @[LZD.scala 43:32]
  wire  _T_346; // @[LZD.scala 39:14]
  wire  _T_347; // @[LZD.scala 39:21]
  wire  _T_348; // @[LZD.scala 39:30]
  wire  _T_349; // @[LZD.scala 39:27]
  wire  _T_350; // @[LZD.scala 39:25]
  wire [1:0] _T_351; // @[Cat.scala 29:58]
  wire [1:0] _T_352; // @[LZD.scala 44:32]
  wire  _T_353; // @[LZD.scala 39:14]
  wire  _T_354; // @[LZD.scala 39:21]
  wire  _T_355; // @[LZD.scala 39:30]
  wire  _T_356; // @[LZD.scala 39:27]
  wire  _T_357; // @[LZD.scala 39:25]
  wire [1:0] _T_358; // @[Cat.scala 29:58]
  wire  _T_359; // @[Shift.scala 12:21]
  wire  _T_360; // @[Shift.scala 12:21]
  wire  _T_361; // @[LZD.scala 49:16]
  wire  _T_362; // @[LZD.scala 49:27]
  wire  _T_363; // @[LZD.scala 49:25]
  wire  _T_364; // @[LZD.scala 49:47]
  wire  _T_365; // @[LZD.scala 49:59]
  wire  _T_366; // @[LZD.scala 49:35]
  wire [2:0] _T_368; // @[Cat.scala 29:58]
  wire [3:0] _T_369; // @[LZD.scala 44:32]
  wire [1:0] _T_370; // @[LZD.scala 43:32]
  wire  _T_371; // @[LZD.scala 39:14]
  wire  _T_372; // @[LZD.scala 39:21]
  wire  _T_373; // @[LZD.scala 39:30]
  wire  _T_374; // @[LZD.scala 39:27]
  wire  _T_375; // @[LZD.scala 39:25]
  wire [1:0] _T_376; // @[Cat.scala 29:58]
  wire [1:0] _T_377; // @[LZD.scala 44:32]
  wire  _T_378; // @[LZD.scala 39:14]
  wire  _T_379; // @[LZD.scala 39:21]
  wire  _T_380; // @[LZD.scala 39:30]
  wire  _T_381; // @[LZD.scala 39:27]
  wire  _T_382; // @[LZD.scala 39:25]
  wire [1:0] _T_383; // @[Cat.scala 29:58]
  wire  _T_384; // @[Shift.scala 12:21]
  wire  _T_385; // @[Shift.scala 12:21]
  wire  _T_386; // @[LZD.scala 49:16]
  wire  _T_387; // @[LZD.scala 49:27]
  wire  _T_388; // @[LZD.scala 49:25]
  wire  _T_389; // @[LZD.scala 49:47]
  wire  _T_390; // @[LZD.scala 49:59]
  wire  _T_391; // @[LZD.scala 49:35]
  wire [2:0] _T_393; // @[Cat.scala 29:58]
  wire  _T_394; // @[Shift.scala 12:21]
  wire  _T_395; // @[Shift.scala 12:21]
  wire  _T_396; // @[LZD.scala 49:16]
  wire  _T_397; // @[LZD.scala 49:27]
  wire  _T_398; // @[LZD.scala 49:25]
  wire [1:0] _T_399; // @[LZD.scala 49:47]
  wire [1:0] _T_400; // @[LZD.scala 49:59]
  wire [1:0] _T_401; // @[LZD.scala 49:35]
  wire [3:0] _T_403; // @[Cat.scala 29:58]
  wire [5:0] _T_404; // @[LZD.scala 44:32]
  wire [3:0] _T_405; // @[LZD.scala 43:32]
  wire [1:0] _T_406; // @[LZD.scala 43:32]
  wire  _T_407; // @[LZD.scala 39:14]
  wire  _T_408; // @[LZD.scala 39:21]
  wire  _T_409; // @[LZD.scala 39:30]
  wire  _T_410; // @[LZD.scala 39:27]
  wire  _T_411; // @[LZD.scala 39:25]
  wire [1:0] _T_412; // @[Cat.scala 29:58]
  wire [1:0] _T_413; // @[LZD.scala 44:32]
  wire  _T_414; // @[LZD.scala 39:14]
  wire  _T_415; // @[LZD.scala 39:21]
  wire  _T_416; // @[LZD.scala 39:30]
  wire  _T_417; // @[LZD.scala 39:27]
  wire  _T_418; // @[LZD.scala 39:25]
  wire [1:0] _T_419; // @[Cat.scala 29:58]
  wire  _T_420; // @[Shift.scala 12:21]
  wire  _T_421; // @[Shift.scala 12:21]
  wire  _T_422; // @[LZD.scala 49:16]
  wire  _T_423; // @[LZD.scala 49:27]
  wire  _T_424; // @[LZD.scala 49:25]
  wire  _T_425; // @[LZD.scala 49:47]
  wire  _T_426; // @[LZD.scala 49:59]
  wire  _T_427; // @[LZD.scala 49:35]
  wire [2:0] _T_429; // @[Cat.scala 29:58]
  wire [1:0] _T_430; // @[LZD.scala 44:32]
  wire  _T_431; // @[LZD.scala 39:14]
  wire  _T_432; // @[LZD.scala 39:21]
  wire  _T_433; // @[LZD.scala 39:30]
  wire  _T_434; // @[LZD.scala 39:27]
  wire  _T_435; // @[LZD.scala 39:25]
  wire [1:0] _T_436; // @[Cat.scala 29:58]
  wire  _T_437; // @[Shift.scala 12:21]
  wire [1:0] _T_439; // @[LZD.scala 55:32]
  wire [1:0] _T_440; // @[LZD.scala 55:20]
  wire [2:0] _T_441; // @[Cat.scala 29:58]
  wire  _T_442; // @[Shift.scala 12:21]
  wire [2:0] _T_444; // @[LZD.scala 55:32]
  wire [2:0] _T_445; // @[LZD.scala 55:20]
  wire [3:0] sumLZD; // @[Cat.scala 29:58]
  wire [4:0] _T_446; // @[Cat.scala 29:58]
  wire [4:0] _T_447; // @[PositAdder.scala 41:38]
  wire [4:0] _T_449; // @[PositAdder.scala 41:45]
  wire [4:0] scaleBias; // @[PositAdder.scala 41:45]
  wire [5:0] _GEN_4; // @[PositAdder.scala 42:32]
  wire [6:0] sumScale; // @[PositAdder.scala 42:32]
  wire  overflow; // @[PositAdder.scala 43:30]
  wire [3:0] normalShift; // @[PositAdder.scala 44:22]
  wire [12:0] _T_450; // @[PositAdder.scala 45:36]
  wire  _T_451; // @[Shift.scala 16:24]
  wire  _T_453; // @[Shift.scala 12:21]
  wire [4:0] _T_454; // @[Shift.scala 64:52]
  wire [12:0] _T_456; // @[Cat.scala 29:58]
  wire [12:0] _T_457; // @[Shift.scala 64:27]
  wire [2:0] _T_458; // @[Shift.scala 66:70]
  wire  _T_459; // @[Shift.scala 12:21]
  wire [8:0] _T_460; // @[Shift.scala 64:52]
  wire [12:0] _T_462; // @[Cat.scala 29:58]
  wire [12:0] _T_463; // @[Shift.scala 64:27]
  wire [1:0] _T_464; // @[Shift.scala 66:70]
  wire  _T_465; // @[Shift.scala 12:21]
  wire [10:0] _T_466; // @[Shift.scala 64:52]
  wire [12:0] _T_468; // @[Cat.scala 29:58]
  wire [12:0] _T_469; // @[Shift.scala 64:27]
  wire  _T_470; // @[Shift.scala 66:70]
  wire [11:0] _T_472; // @[Shift.scala 64:52]
  wire [12:0] _T_473; // @[Cat.scala 29:58]
  wire [12:0] _T_474; // @[Shift.scala 64:27]
  wire [12:0] shiftSig; // @[Shift.scala 16:10]
  wire [6:0] _T_475; // @[PositAdder.scala 50:24]
  wire [8:0] decS_fraction; // @[PositAdder.scala 51:34]
  wire  decS_isNaR; // @[PositAdder.scala 52:32]
  wire  _T_478; // @[PositAdder.scala 53:33]
  wire  _T_479; // @[PositAdder.scala 53:21]
  wire  _T_480; // @[PositAdder.scala 53:52]
  wire  decS_isZero; // @[PositAdder.scala 53:37]
  wire [1:0] _T_482; // @[PositAdder.scala 54:33]
  wire  _T_483; // @[PositAdder.scala 54:49]
  wire  _T_484; // @[PositAdder.scala 54:63]
  wire  _T_485; // @[PositAdder.scala 54:53]
  wire [5:0] _GEN_5; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  wire [5:0] decS_scale; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  wire  _T_488; // @[convert.scala 46:61]
  wire  _T_489; // @[convert.scala 46:52]
  wire  _T_491; // @[convert.scala 46:42]
  wire [4:0] _T_492; // @[convert.scala 48:34]
  wire  _T_493; // @[convert.scala 49:36]
  wire [4:0] _T_495; // @[convert.scala 50:36]
  wire [4:0] _T_496; // @[convert.scala 50:36]
  wire [4:0] _T_497; // @[convert.scala 50:28]
  wire  _T_498; // @[convert.scala 51:31]
  wire  _T_499; // @[convert.scala 52:43]
  wire [14:0] _T_503; // @[Cat.scala 29:58]
  wire [4:0] _T_504; // @[Shift.scala 39:17]
  wire  _T_505; // @[Shift.scala 39:24]
  wire [3:0] _T_506; // @[Shift.scala 40:44]
  wire [6:0] _T_507; // @[Shift.scala 90:30]
  wire [7:0] _T_508; // @[Shift.scala 90:48]
  wire  _T_509; // @[Shift.scala 90:57]
  wire [6:0] _GEN_6; // @[Shift.scala 90:39]
  wire [6:0] _T_510; // @[Shift.scala 90:39]
  wire  _T_511; // @[Shift.scala 12:21]
  wire  _T_512; // @[Shift.scala 12:21]
  wire [7:0] _T_514; // @[Bitwise.scala 71:12]
  wire [14:0] _T_515; // @[Cat.scala 29:58]
  wire [14:0] _T_516; // @[Shift.scala 91:22]
  wire [2:0] _T_517; // @[Shift.scala 92:77]
  wire [10:0] _T_518; // @[Shift.scala 90:30]
  wire [3:0] _T_519; // @[Shift.scala 90:48]
  wire  _T_520; // @[Shift.scala 90:57]
  wire [10:0] _GEN_7; // @[Shift.scala 90:39]
  wire [10:0] _T_521; // @[Shift.scala 90:39]
  wire  _T_522; // @[Shift.scala 12:21]
  wire  _T_523; // @[Shift.scala 12:21]
  wire [3:0] _T_525; // @[Bitwise.scala 71:12]
  wire [14:0] _T_526; // @[Cat.scala 29:58]
  wire [14:0] _T_527; // @[Shift.scala 91:22]
  wire [1:0] _T_528; // @[Shift.scala 92:77]
  wire [12:0] _T_529; // @[Shift.scala 90:30]
  wire [1:0] _T_530; // @[Shift.scala 90:48]
  wire  _T_531; // @[Shift.scala 90:57]
  wire [12:0] _GEN_8; // @[Shift.scala 90:39]
  wire [12:0] _T_532; // @[Shift.scala 90:39]
  wire  _T_533; // @[Shift.scala 12:21]
  wire  _T_534; // @[Shift.scala 12:21]
  wire [1:0] _T_536; // @[Bitwise.scala 71:12]
  wire [14:0] _T_537; // @[Cat.scala 29:58]
  wire [14:0] _T_538; // @[Shift.scala 91:22]
  wire  _T_539; // @[Shift.scala 92:77]
  wire [13:0] _T_540; // @[Shift.scala 90:30]
  wire  _T_541; // @[Shift.scala 90:48]
  wire [13:0] _GEN_9; // @[Shift.scala 90:39]
  wire [13:0] _T_543; // @[Shift.scala 90:39]
  wire  _T_545; // @[Shift.scala 12:21]
  wire [14:0] _T_546; // @[Cat.scala 29:58]
  wire [14:0] _T_547; // @[Shift.scala 91:22]
  wire [14:0] _T_550; // @[Bitwise.scala 71:12]
  wire [14:0] _T_551; // @[Shift.scala 39:10]
  wire  _T_552; // @[convert.scala 55:31]
  wire  _T_553; // @[convert.scala 56:31]
  wire  _T_554; // @[convert.scala 57:31]
  wire  _T_555; // @[convert.scala 58:31]
  wire [11:0] _T_556; // @[convert.scala 59:69]
  wire  _T_557; // @[convert.scala 59:81]
  wire  _T_558; // @[convert.scala 59:50]
  wire  _T_560; // @[convert.scala 60:81]
  wire  _T_561; // @[convert.scala 61:44]
  wire  _T_562; // @[convert.scala 61:52]
  wire  _T_563; // @[convert.scala 61:36]
  wire  _T_564; // @[convert.scala 62:63]
  wire  _T_565; // @[convert.scala 62:103]
  wire  _T_566; // @[convert.scala 62:60]
  wire [11:0] _GEN_10; // @[convert.scala 63:56]
  wire [11:0] _T_569; // @[convert.scala 63:56]
  wire [12:0] _T_570; // @[Cat.scala 29:58]
  wire [12:0] _T_572; // @[Mux.scala 87:16]
  assign _T_1 = io_A[12]; // @[convert.scala 18:24]
  assign _T_2 = io_A[11]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[11:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[10:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[10:3]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[2:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68[2:1]; // @[LZD.scala 43:32]
  assign _T_70 = _T_69 != 2'h0; // @[LZD.scala 39:14]
  assign _T_71 = _T_69[1]; // @[LZD.scala 39:21]
  assign _T_72 = _T_69[0]; // @[LZD.scala 39:30]
  assign _T_73 = ~ _T_72; // @[LZD.scala 39:27]
  assign _T_74 = _T_71 | _T_73; // @[LZD.scala 39:25]
  assign _T_75 = {_T_70,_T_74}; // @[Cat.scala 29:58]
  assign _T_76 = _T_68[0:0]; // @[LZD.scala 44:32]
  assign _T_78 = _T_75[1]; // @[Shift.scala 12:21]
  assign _T_80 = _T_75[0:0]; // @[LZD.scala 55:32]
  assign _T_81 = _T_78 ? _T_80 : _T_76; // @[LZD.scala 55:20]
  assign _T_83 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_85 = {1'h1,_T_78,_T_81}; // @[Cat.scala 29:58]
  assign _T_86 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_87 = _T_83 ? _T_86 : _T_85; // @[LZD.scala 55:20]
  assign _T_88 = {_T_83,_T_87}; // @[Cat.scala 29:58]
  assign _T_89 = ~ _T_88; // @[convert.scala 21:22]
  assign _T_90 = io_A[9:0]; // @[convert.scala 22:36]
  assign _T_91 = _T_89 < 4'ha; // @[Shift.scala 16:24]
  assign _T_93 = _T_89[3]; // @[Shift.scala 12:21]
  assign _T_94 = _T_90[1:0]; // @[Shift.scala 64:52]
  assign _T_96 = {_T_94,8'h0}; // @[Cat.scala 29:58]
  assign _T_97 = _T_93 ? _T_96 : _T_90; // @[Shift.scala 64:27]
  assign _T_98 = _T_89[2:0]; // @[Shift.scala 66:70]
  assign _T_99 = _T_98[2]; // @[Shift.scala 12:21]
  assign _T_100 = _T_97[5:0]; // @[Shift.scala 64:52]
  assign _T_102 = {_T_100,4'h0}; // @[Cat.scala 29:58]
  assign _T_103 = _T_99 ? _T_102 : _T_97; // @[Shift.scala 64:27]
  assign _T_104 = _T_98[1:0]; // @[Shift.scala 66:70]
  assign _T_105 = _T_104[1]; // @[Shift.scala 12:21]
  assign _T_106 = _T_103[7:0]; // @[Shift.scala 64:52]
  assign _T_108 = {_T_106,2'h0}; // @[Cat.scala 29:58]
  assign _T_109 = _T_105 ? _T_108 : _T_103; // @[Shift.scala 64:27]
  assign _T_110 = _T_104[0:0]; // @[Shift.scala 66:70]
  assign _T_112 = _T_109[8:0]; // @[Shift.scala 64:52]
  assign _T_113 = {_T_112,1'h0}; // @[Cat.scala 29:58]
  assign _T_114 = _T_110 ? _T_113 : _T_109; // @[Shift.scala 64:27]
  assign _T_115 = _T_91 ? _T_114 : 10'h0; // @[Shift.scala 16:10]
  assign _T_116 = _T_115[9:9]; // @[convert.scala 23:34]
  assign decA_fraction = _T_115[8:0]; // @[convert.scala 24:34]
  assign _T_118 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_120 = _T_3 ? _T_89 : _T_88; // @[convert.scala 25:42]
  assign _T_123 = ~ _T_116; // @[convert.scala 26:67]
  assign _T_124 = _T_1 ? _T_123 : _T_116; // @[convert.scala 26:51]
  assign _T_125 = {_T_118,_T_120,_T_124}; // @[Cat.scala 29:58]
  assign _T_127 = io_A[11:0]; // @[convert.scala 29:56]
  assign _T_128 = _T_127 != 12'h0; // @[convert.scala 29:60]
  assign _T_129 = ~ _T_128; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_129; // @[convert.scala 29:39]
  assign _T_132 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_132 & _T_129; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_125); // @[convert.scala 32:24]
  assign _T_141 = io_B[12]; // @[convert.scala 18:24]
  assign _T_142 = io_B[11]; // @[convert.scala 18:40]
  assign _T_143 = _T_141 ^ _T_142; // @[convert.scala 18:36]
  assign _T_144 = io_B[11:1]; // @[convert.scala 19:24]
  assign _T_145 = io_B[10:0]; // @[convert.scala 19:43]
  assign _T_146 = _T_144 ^ _T_145; // @[convert.scala 19:39]
  assign _T_147 = _T_146[10:3]; // @[LZD.scala 43:32]
  assign _T_148 = _T_147[7:4]; // @[LZD.scala 43:32]
  assign _T_149 = _T_148[3:2]; // @[LZD.scala 43:32]
  assign _T_150 = _T_149 != 2'h0; // @[LZD.scala 39:14]
  assign _T_151 = _T_149[1]; // @[LZD.scala 39:21]
  assign _T_152 = _T_149[0]; // @[LZD.scala 39:30]
  assign _T_153 = ~ _T_152; // @[LZD.scala 39:27]
  assign _T_154 = _T_151 | _T_153; // @[LZD.scala 39:25]
  assign _T_155 = {_T_150,_T_154}; // @[Cat.scala 29:58]
  assign _T_156 = _T_148[1:0]; // @[LZD.scala 44:32]
  assign _T_157 = _T_156 != 2'h0; // @[LZD.scala 39:14]
  assign _T_158 = _T_156[1]; // @[LZD.scala 39:21]
  assign _T_159 = _T_156[0]; // @[LZD.scala 39:30]
  assign _T_160 = ~ _T_159; // @[LZD.scala 39:27]
  assign _T_161 = _T_158 | _T_160; // @[LZD.scala 39:25]
  assign _T_162 = {_T_157,_T_161}; // @[Cat.scala 29:58]
  assign _T_163 = _T_155[1]; // @[Shift.scala 12:21]
  assign _T_164 = _T_162[1]; // @[Shift.scala 12:21]
  assign _T_165 = _T_163 | _T_164; // @[LZD.scala 49:16]
  assign _T_166 = ~ _T_164; // @[LZD.scala 49:27]
  assign _T_167 = _T_163 | _T_166; // @[LZD.scala 49:25]
  assign _T_168 = _T_155[0:0]; // @[LZD.scala 49:47]
  assign _T_169 = _T_162[0:0]; // @[LZD.scala 49:59]
  assign _T_170 = _T_163 ? _T_168 : _T_169; // @[LZD.scala 49:35]
  assign _T_172 = {_T_165,_T_167,_T_170}; // @[Cat.scala 29:58]
  assign _T_173 = _T_147[3:0]; // @[LZD.scala 44:32]
  assign _T_174 = _T_173[3:2]; // @[LZD.scala 43:32]
  assign _T_175 = _T_174 != 2'h0; // @[LZD.scala 39:14]
  assign _T_176 = _T_174[1]; // @[LZD.scala 39:21]
  assign _T_177 = _T_174[0]; // @[LZD.scala 39:30]
  assign _T_178 = ~ _T_177; // @[LZD.scala 39:27]
  assign _T_179 = _T_176 | _T_178; // @[LZD.scala 39:25]
  assign _T_180 = {_T_175,_T_179}; // @[Cat.scala 29:58]
  assign _T_181 = _T_173[1:0]; // @[LZD.scala 44:32]
  assign _T_182 = _T_181 != 2'h0; // @[LZD.scala 39:14]
  assign _T_183 = _T_181[1]; // @[LZD.scala 39:21]
  assign _T_184 = _T_181[0]; // @[LZD.scala 39:30]
  assign _T_185 = ~ _T_184; // @[LZD.scala 39:27]
  assign _T_186 = _T_183 | _T_185; // @[LZD.scala 39:25]
  assign _T_187 = {_T_182,_T_186}; // @[Cat.scala 29:58]
  assign _T_188 = _T_180[1]; // @[Shift.scala 12:21]
  assign _T_189 = _T_187[1]; // @[Shift.scala 12:21]
  assign _T_190 = _T_188 | _T_189; // @[LZD.scala 49:16]
  assign _T_191 = ~ _T_189; // @[LZD.scala 49:27]
  assign _T_192 = _T_188 | _T_191; // @[LZD.scala 49:25]
  assign _T_193 = _T_180[0:0]; // @[LZD.scala 49:47]
  assign _T_194 = _T_187[0:0]; // @[LZD.scala 49:59]
  assign _T_195 = _T_188 ? _T_193 : _T_194; // @[LZD.scala 49:35]
  assign _T_197 = {_T_190,_T_192,_T_195}; // @[Cat.scala 29:58]
  assign _T_198 = _T_172[2]; // @[Shift.scala 12:21]
  assign _T_199 = _T_197[2]; // @[Shift.scala 12:21]
  assign _T_200 = _T_198 | _T_199; // @[LZD.scala 49:16]
  assign _T_201 = ~ _T_199; // @[LZD.scala 49:27]
  assign _T_202 = _T_198 | _T_201; // @[LZD.scala 49:25]
  assign _T_203 = _T_172[1:0]; // @[LZD.scala 49:47]
  assign _T_204 = _T_197[1:0]; // @[LZD.scala 49:59]
  assign _T_205 = _T_198 ? _T_203 : _T_204; // @[LZD.scala 49:35]
  assign _T_207 = {_T_200,_T_202,_T_205}; // @[Cat.scala 29:58]
  assign _T_208 = _T_146[2:0]; // @[LZD.scala 44:32]
  assign _T_209 = _T_208[2:1]; // @[LZD.scala 43:32]
  assign _T_210 = _T_209 != 2'h0; // @[LZD.scala 39:14]
  assign _T_211 = _T_209[1]; // @[LZD.scala 39:21]
  assign _T_212 = _T_209[0]; // @[LZD.scala 39:30]
  assign _T_213 = ~ _T_212; // @[LZD.scala 39:27]
  assign _T_214 = _T_211 | _T_213; // @[LZD.scala 39:25]
  assign _T_215 = {_T_210,_T_214}; // @[Cat.scala 29:58]
  assign _T_216 = _T_208[0:0]; // @[LZD.scala 44:32]
  assign _T_218 = _T_215[1]; // @[Shift.scala 12:21]
  assign _T_220 = _T_215[0:0]; // @[LZD.scala 55:32]
  assign _T_221 = _T_218 ? _T_220 : _T_216; // @[LZD.scala 55:20]
  assign _T_223 = _T_207[3]; // @[Shift.scala 12:21]
  assign _T_225 = {1'h1,_T_218,_T_221}; // @[Cat.scala 29:58]
  assign _T_226 = _T_207[2:0]; // @[LZD.scala 55:32]
  assign _T_227 = _T_223 ? _T_226 : _T_225; // @[LZD.scala 55:20]
  assign _T_228 = {_T_223,_T_227}; // @[Cat.scala 29:58]
  assign _T_229 = ~ _T_228; // @[convert.scala 21:22]
  assign _T_230 = io_B[9:0]; // @[convert.scala 22:36]
  assign _T_231 = _T_229 < 4'ha; // @[Shift.scala 16:24]
  assign _T_233 = _T_229[3]; // @[Shift.scala 12:21]
  assign _T_234 = _T_230[1:0]; // @[Shift.scala 64:52]
  assign _T_236 = {_T_234,8'h0}; // @[Cat.scala 29:58]
  assign _T_237 = _T_233 ? _T_236 : _T_230; // @[Shift.scala 64:27]
  assign _T_238 = _T_229[2:0]; // @[Shift.scala 66:70]
  assign _T_239 = _T_238[2]; // @[Shift.scala 12:21]
  assign _T_240 = _T_237[5:0]; // @[Shift.scala 64:52]
  assign _T_242 = {_T_240,4'h0}; // @[Cat.scala 29:58]
  assign _T_243 = _T_239 ? _T_242 : _T_237; // @[Shift.scala 64:27]
  assign _T_244 = _T_238[1:0]; // @[Shift.scala 66:70]
  assign _T_245 = _T_244[1]; // @[Shift.scala 12:21]
  assign _T_246 = _T_243[7:0]; // @[Shift.scala 64:52]
  assign _T_248 = {_T_246,2'h0}; // @[Cat.scala 29:58]
  assign _T_249 = _T_245 ? _T_248 : _T_243; // @[Shift.scala 64:27]
  assign _T_250 = _T_244[0:0]; // @[Shift.scala 66:70]
  assign _T_252 = _T_249[8:0]; // @[Shift.scala 64:52]
  assign _T_253 = {_T_252,1'h0}; // @[Cat.scala 29:58]
  assign _T_254 = _T_250 ? _T_253 : _T_249; // @[Shift.scala 64:27]
  assign _T_255 = _T_231 ? _T_254 : 10'h0; // @[Shift.scala 16:10]
  assign _T_256 = _T_255[9:9]; // @[convert.scala 23:34]
  assign decB_fraction = _T_255[8:0]; // @[convert.scala 24:34]
  assign _T_258 = _T_143 == 1'h0; // @[convert.scala 25:26]
  assign _T_260 = _T_143 ? _T_229 : _T_228; // @[convert.scala 25:42]
  assign _T_263 = ~ _T_256; // @[convert.scala 26:67]
  assign _T_264 = _T_141 ? _T_263 : _T_256; // @[convert.scala 26:51]
  assign _T_265 = {_T_258,_T_260,_T_264}; // @[Cat.scala 29:58]
  assign _T_267 = io_B[11:0]; // @[convert.scala 29:56]
  assign _T_268 = _T_267 != 12'h0; // @[convert.scala 29:60]
  assign _T_269 = ~ _T_268; // @[convert.scala 29:41]
  assign decB_isNaR = _T_141 & _T_269; // @[convert.scala 29:39]
  assign _T_272 = _T_141 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_272 & _T_269; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_265); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[PositAdder.scala 24:32]
  assign greaterSign = aGTb ? _T_1 : _T_141; // @[PositAdder.scala 25:24]
  assign smallerSign = aGTb ? _T_141 : _T_1; // @[PositAdder.scala 26:24]
  assign greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[PositAdder.scala 27:24]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[PositAdder.scala 28:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[PositAdder.scala 29:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[PositAdder.scala 30:24]
  assign _T_281 = $signed(greaterExp) - $signed(smallerExp); // @[PositAdder.scala 31:32]
  assign scale_diff = $signed(_T_281); // @[PositAdder.scala 31:32]
  assign _T_282 = ~ greaterSign; // @[PositAdder.scala 32:38]
  assign greaterSig = {greaterSign,_T_282,greaterFrac}; // @[Cat.scala 29:58]
  assign _T_284 = ~ smallerSign; // @[PositAdder.scala 33:38]
  assign _T_287 = {smallerSign,_T_284,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_288 = $unsigned(scale_diff); // @[PositAdder.scala 34:68]
  assign _T_289 = _T_288 < 6'he; // @[Shift.scala 39:24]
  assign _T_290 = _T_288[3:0]; // @[Shift.scala 40:44]
  assign _T_291 = _T_287[13:8]; // @[Shift.scala 90:30]
  assign _T_292 = _T_287[7:0]; // @[Shift.scala 90:48]
  assign _T_293 = _T_292 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{5'd0}, _T_293}; // @[Shift.scala 90:39]
  assign _T_294 = _T_291 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_295 = _T_290[3]; // @[Shift.scala 12:21]
  assign _T_296 = _T_287[13]; // @[Shift.scala 12:21]
  assign _T_298 = _T_296 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_299 = {_T_298,_T_294}; // @[Cat.scala 29:58]
  assign _T_300 = _T_295 ? _T_299 : _T_287; // @[Shift.scala 91:22]
  assign _T_301 = _T_290[2:0]; // @[Shift.scala 92:77]
  assign _T_302 = _T_300[13:4]; // @[Shift.scala 90:30]
  assign _T_303 = _T_300[3:0]; // @[Shift.scala 90:48]
  assign _T_304 = _T_303 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{9'd0}, _T_304}; // @[Shift.scala 90:39]
  assign _T_305 = _T_302 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_306 = _T_301[2]; // @[Shift.scala 12:21]
  assign _T_307 = _T_300[13]; // @[Shift.scala 12:21]
  assign _T_309 = _T_307 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_310 = {_T_309,_T_305}; // @[Cat.scala 29:58]
  assign _T_311 = _T_306 ? _T_310 : _T_300; // @[Shift.scala 91:22]
  assign _T_312 = _T_301[1:0]; // @[Shift.scala 92:77]
  assign _T_313 = _T_311[13:2]; // @[Shift.scala 90:30]
  assign _T_314 = _T_311[1:0]; // @[Shift.scala 90:48]
  assign _T_315 = _T_314 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{11'd0}, _T_315}; // @[Shift.scala 90:39]
  assign _T_316 = _T_313 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_317 = _T_312[1]; // @[Shift.scala 12:21]
  assign _T_318 = _T_311[13]; // @[Shift.scala 12:21]
  assign _T_320 = _T_318 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_321 = {_T_320,_T_316}; // @[Cat.scala 29:58]
  assign _T_322 = _T_317 ? _T_321 : _T_311; // @[Shift.scala 91:22]
  assign _T_323 = _T_312[0:0]; // @[Shift.scala 92:77]
  assign _T_324 = _T_322[13:1]; // @[Shift.scala 90:30]
  assign _T_325 = _T_322[0:0]; // @[Shift.scala 90:48]
  assign _GEN_3 = {{12'd0}, _T_325}; // @[Shift.scala 90:39]
  assign _T_327 = _T_324 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_329 = _T_322[13]; // @[Shift.scala 12:21]
  assign _T_330 = {_T_329,_T_327}; // @[Cat.scala 29:58]
  assign _T_331 = _T_323 ? _T_330 : _T_322; // @[Shift.scala 91:22]
  assign _T_334 = _T_296 ? 14'h3fff : 14'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_289 ? _T_331 : _T_334; // @[Shift.scala 39:10]
  assign _T_335 = smallerSig[13:3]; // @[PositAdder.scala 35:45]
  assign rawSumSig = greaterSig + _T_335; // @[PositAdder.scala 35:32]
  assign _T_336 = _T_1 ^ _T_141; // @[PositAdder.scala 36:31]
  assign _T_337 = rawSumSig[11:11]; // @[PositAdder.scala 36:59]
  assign sumSign = _T_336 ^ _T_337; // @[PositAdder.scala 36:43]
  assign _T_338 = greaterSig + _T_335; // @[PositAdder.scala 37:48]
  assign _T_339 = smallerSig[2:0]; // @[PositAdder.scala 37:63]
  assign signSumSig = {sumSign,_T_338,_T_339}; // @[Cat.scala 29:58]
  assign _T_341 = signSumSig[14:1]; // @[PositAdder.scala 39:31]
  assign _T_342 = signSumSig[13:0]; // @[PositAdder.scala 39:66]
  assign sumXor = _T_341 ^ _T_342; // @[PositAdder.scala 39:49]
  assign _T_343 = sumXor[13:6]; // @[LZD.scala 43:32]
  assign _T_344 = _T_343[7:4]; // @[LZD.scala 43:32]
  assign _T_345 = _T_344[3:2]; // @[LZD.scala 43:32]
  assign _T_346 = _T_345 != 2'h0; // @[LZD.scala 39:14]
  assign _T_347 = _T_345[1]; // @[LZD.scala 39:21]
  assign _T_348 = _T_345[0]; // @[LZD.scala 39:30]
  assign _T_349 = ~ _T_348; // @[LZD.scala 39:27]
  assign _T_350 = _T_347 | _T_349; // @[LZD.scala 39:25]
  assign _T_351 = {_T_346,_T_350}; // @[Cat.scala 29:58]
  assign _T_352 = _T_344[1:0]; // @[LZD.scala 44:32]
  assign _T_353 = _T_352 != 2'h0; // @[LZD.scala 39:14]
  assign _T_354 = _T_352[1]; // @[LZD.scala 39:21]
  assign _T_355 = _T_352[0]; // @[LZD.scala 39:30]
  assign _T_356 = ~ _T_355; // @[LZD.scala 39:27]
  assign _T_357 = _T_354 | _T_356; // @[LZD.scala 39:25]
  assign _T_358 = {_T_353,_T_357}; // @[Cat.scala 29:58]
  assign _T_359 = _T_351[1]; // @[Shift.scala 12:21]
  assign _T_360 = _T_358[1]; // @[Shift.scala 12:21]
  assign _T_361 = _T_359 | _T_360; // @[LZD.scala 49:16]
  assign _T_362 = ~ _T_360; // @[LZD.scala 49:27]
  assign _T_363 = _T_359 | _T_362; // @[LZD.scala 49:25]
  assign _T_364 = _T_351[0:0]; // @[LZD.scala 49:47]
  assign _T_365 = _T_358[0:0]; // @[LZD.scala 49:59]
  assign _T_366 = _T_359 ? _T_364 : _T_365; // @[LZD.scala 49:35]
  assign _T_368 = {_T_361,_T_363,_T_366}; // @[Cat.scala 29:58]
  assign _T_369 = _T_343[3:0]; // @[LZD.scala 44:32]
  assign _T_370 = _T_369[3:2]; // @[LZD.scala 43:32]
  assign _T_371 = _T_370 != 2'h0; // @[LZD.scala 39:14]
  assign _T_372 = _T_370[1]; // @[LZD.scala 39:21]
  assign _T_373 = _T_370[0]; // @[LZD.scala 39:30]
  assign _T_374 = ~ _T_373; // @[LZD.scala 39:27]
  assign _T_375 = _T_372 | _T_374; // @[LZD.scala 39:25]
  assign _T_376 = {_T_371,_T_375}; // @[Cat.scala 29:58]
  assign _T_377 = _T_369[1:0]; // @[LZD.scala 44:32]
  assign _T_378 = _T_377 != 2'h0; // @[LZD.scala 39:14]
  assign _T_379 = _T_377[1]; // @[LZD.scala 39:21]
  assign _T_380 = _T_377[0]; // @[LZD.scala 39:30]
  assign _T_381 = ~ _T_380; // @[LZD.scala 39:27]
  assign _T_382 = _T_379 | _T_381; // @[LZD.scala 39:25]
  assign _T_383 = {_T_378,_T_382}; // @[Cat.scala 29:58]
  assign _T_384 = _T_376[1]; // @[Shift.scala 12:21]
  assign _T_385 = _T_383[1]; // @[Shift.scala 12:21]
  assign _T_386 = _T_384 | _T_385; // @[LZD.scala 49:16]
  assign _T_387 = ~ _T_385; // @[LZD.scala 49:27]
  assign _T_388 = _T_384 | _T_387; // @[LZD.scala 49:25]
  assign _T_389 = _T_376[0:0]; // @[LZD.scala 49:47]
  assign _T_390 = _T_383[0:0]; // @[LZD.scala 49:59]
  assign _T_391 = _T_384 ? _T_389 : _T_390; // @[LZD.scala 49:35]
  assign _T_393 = {_T_386,_T_388,_T_391}; // @[Cat.scala 29:58]
  assign _T_394 = _T_368[2]; // @[Shift.scala 12:21]
  assign _T_395 = _T_393[2]; // @[Shift.scala 12:21]
  assign _T_396 = _T_394 | _T_395; // @[LZD.scala 49:16]
  assign _T_397 = ~ _T_395; // @[LZD.scala 49:27]
  assign _T_398 = _T_394 | _T_397; // @[LZD.scala 49:25]
  assign _T_399 = _T_368[1:0]; // @[LZD.scala 49:47]
  assign _T_400 = _T_393[1:0]; // @[LZD.scala 49:59]
  assign _T_401 = _T_394 ? _T_399 : _T_400; // @[LZD.scala 49:35]
  assign _T_403 = {_T_396,_T_398,_T_401}; // @[Cat.scala 29:58]
  assign _T_404 = sumXor[5:0]; // @[LZD.scala 44:32]
  assign _T_405 = _T_404[5:2]; // @[LZD.scala 43:32]
  assign _T_406 = _T_405[3:2]; // @[LZD.scala 43:32]
  assign _T_407 = _T_406 != 2'h0; // @[LZD.scala 39:14]
  assign _T_408 = _T_406[1]; // @[LZD.scala 39:21]
  assign _T_409 = _T_406[0]; // @[LZD.scala 39:30]
  assign _T_410 = ~ _T_409; // @[LZD.scala 39:27]
  assign _T_411 = _T_408 | _T_410; // @[LZD.scala 39:25]
  assign _T_412 = {_T_407,_T_411}; // @[Cat.scala 29:58]
  assign _T_413 = _T_405[1:0]; // @[LZD.scala 44:32]
  assign _T_414 = _T_413 != 2'h0; // @[LZD.scala 39:14]
  assign _T_415 = _T_413[1]; // @[LZD.scala 39:21]
  assign _T_416 = _T_413[0]; // @[LZD.scala 39:30]
  assign _T_417 = ~ _T_416; // @[LZD.scala 39:27]
  assign _T_418 = _T_415 | _T_417; // @[LZD.scala 39:25]
  assign _T_419 = {_T_414,_T_418}; // @[Cat.scala 29:58]
  assign _T_420 = _T_412[1]; // @[Shift.scala 12:21]
  assign _T_421 = _T_419[1]; // @[Shift.scala 12:21]
  assign _T_422 = _T_420 | _T_421; // @[LZD.scala 49:16]
  assign _T_423 = ~ _T_421; // @[LZD.scala 49:27]
  assign _T_424 = _T_420 | _T_423; // @[LZD.scala 49:25]
  assign _T_425 = _T_412[0:0]; // @[LZD.scala 49:47]
  assign _T_426 = _T_419[0:0]; // @[LZD.scala 49:59]
  assign _T_427 = _T_420 ? _T_425 : _T_426; // @[LZD.scala 49:35]
  assign _T_429 = {_T_422,_T_424,_T_427}; // @[Cat.scala 29:58]
  assign _T_430 = _T_404[1:0]; // @[LZD.scala 44:32]
  assign _T_431 = _T_430 != 2'h0; // @[LZD.scala 39:14]
  assign _T_432 = _T_430[1]; // @[LZD.scala 39:21]
  assign _T_433 = _T_430[0]; // @[LZD.scala 39:30]
  assign _T_434 = ~ _T_433; // @[LZD.scala 39:27]
  assign _T_435 = _T_432 | _T_434; // @[LZD.scala 39:25]
  assign _T_436 = {_T_431,_T_435}; // @[Cat.scala 29:58]
  assign _T_437 = _T_429[2]; // @[Shift.scala 12:21]
  assign _T_439 = _T_429[1:0]; // @[LZD.scala 55:32]
  assign _T_440 = _T_437 ? _T_439 : _T_436; // @[LZD.scala 55:20]
  assign _T_441 = {_T_437,_T_440}; // @[Cat.scala 29:58]
  assign _T_442 = _T_403[3]; // @[Shift.scala 12:21]
  assign _T_444 = _T_403[2:0]; // @[LZD.scala 55:32]
  assign _T_445 = _T_442 ? _T_444 : _T_441; // @[LZD.scala 55:20]
  assign sumLZD = {_T_442,_T_445}; // @[Cat.scala 29:58]
  assign _T_446 = {1'h1,_T_442,_T_445}; // @[Cat.scala 29:58]
  assign _T_447 = $signed(_T_446); // @[PositAdder.scala 41:38]
  assign _T_449 = $signed(_T_447) + $signed(5'sh2); // @[PositAdder.scala 41:45]
  assign scaleBias = $signed(_T_449); // @[PositAdder.scala 41:45]
  assign _GEN_4 = {{1{scaleBias[4]}},scaleBias}; // @[PositAdder.scala 42:32]
  assign sumScale = $signed(greaterExp) + $signed(_GEN_4); // @[PositAdder.scala 42:32]
  assign overflow = $signed(sumScale) > $signed(7'sh16); // @[PositAdder.scala 43:30]
  assign normalShift = ~ sumLZD; // @[PositAdder.scala 44:22]
  assign _T_450 = signSumSig[12:0]; // @[PositAdder.scala 45:36]
  assign _T_451 = normalShift < 4'hd; // @[Shift.scala 16:24]
  assign _T_453 = normalShift[3]; // @[Shift.scala 12:21]
  assign _T_454 = _T_450[4:0]; // @[Shift.scala 64:52]
  assign _T_456 = {_T_454,8'h0}; // @[Cat.scala 29:58]
  assign _T_457 = _T_453 ? _T_456 : _T_450; // @[Shift.scala 64:27]
  assign _T_458 = normalShift[2:0]; // @[Shift.scala 66:70]
  assign _T_459 = _T_458[2]; // @[Shift.scala 12:21]
  assign _T_460 = _T_457[8:0]; // @[Shift.scala 64:52]
  assign _T_462 = {_T_460,4'h0}; // @[Cat.scala 29:58]
  assign _T_463 = _T_459 ? _T_462 : _T_457; // @[Shift.scala 64:27]
  assign _T_464 = _T_458[1:0]; // @[Shift.scala 66:70]
  assign _T_465 = _T_464[1]; // @[Shift.scala 12:21]
  assign _T_466 = _T_463[10:0]; // @[Shift.scala 64:52]
  assign _T_468 = {_T_466,2'h0}; // @[Cat.scala 29:58]
  assign _T_469 = _T_465 ? _T_468 : _T_463; // @[Shift.scala 64:27]
  assign _T_470 = _T_464[0:0]; // @[Shift.scala 66:70]
  assign _T_472 = _T_469[11:0]; // @[Shift.scala 64:52]
  assign _T_473 = {_T_472,1'h0}; // @[Cat.scala 29:58]
  assign _T_474 = _T_470 ? _T_473 : _T_469; // @[Shift.scala 64:27]
  assign shiftSig = _T_451 ? _T_474 : 13'h0; // @[Shift.scala 16:10]
  assign _T_475 = overflow ? $signed(7'sh16) : $signed(sumScale); // @[PositAdder.scala 50:24]
  assign decS_fraction = shiftSig[12:4]; // @[PositAdder.scala 51:34]
  assign decS_isNaR = decA_isNaR | decB_isNaR; // @[PositAdder.scala 52:32]
  assign _T_478 = signSumSig != 15'h0; // @[PositAdder.scala 53:33]
  assign _T_479 = ~ _T_478; // @[PositAdder.scala 53:21]
  assign _T_480 = decA_isZero & decB_isZero; // @[PositAdder.scala 53:52]
  assign decS_isZero = _T_479 | _T_480; // @[PositAdder.scala 53:37]
  assign _T_482 = shiftSig[3:2]; // @[PositAdder.scala 54:33]
  assign _T_483 = shiftSig[1]; // @[PositAdder.scala 54:49]
  assign _T_484 = shiftSig[0]; // @[PositAdder.scala 54:63]
  assign _T_485 = _T_483 | _T_484; // @[PositAdder.scala 54:53]
  assign _GEN_5 = _T_475[5:0]; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  assign decS_scale = $signed(_GEN_5); // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  assign _T_488 = decS_scale[0]; // @[convert.scala 46:61]
  assign _T_489 = ~ _T_488; // @[convert.scala 46:52]
  assign _T_491 = sumSign ? _T_489 : _T_488; // @[convert.scala 46:42]
  assign _T_492 = decS_scale[5:1]; // @[convert.scala 48:34]
  assign _T_493 = _T_492[4:4]; // @[convert.scala 49:36]
  assign _T_495 = ~ _T_492; // @[convert.scala 50:36]
  assign _T_496 = $signed(_T_495); // @[convert.scala 50:36]
  assign _T_497 = _T_493 ? $signed(_T_496) : $signed(_T_492); // @[convert.scala 50:28]
  assign _T_498 = _T_493 ^ sumSign; // @[convert.scala 51:31]
  assign _T_499 = ~ _T_498; // @[convert.scala 52:43]
  assign _T_503 = {_T_499,_T_498,_T_491,decS_fraction,_T_482,_T_485}; // @[Cat.scala 29:58]
  assign _T_504 = $unsigned(_T_497); // @[Shift.scala 39:17]
  assign _T_505 = _T_504 < 5'hf; // @[Shift.scala 39:24]
  assign _T_506 = _T_497[3:0]; // @[Shift.scala 40:44]
  assign _T_507 = _T_503[14:8]; // @[Shift.scala 90:30]
  assign _T_508 = _T_503[7:0]; // @[Shift.scala 90:48]
  assign _T_509 = _T_508 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{6'd0}, _T_509}; // @[Shift.scala 90:39]
  assign _T_510 = _T_507 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_511 = _T_506[3]; // @[Shift.scala 12:21]
  assign _T_512 = _T_503[14]; // @[Shift.scala 12:21]
  assign _T_514 = _T_512 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_515 = {_T_514,_T_510}; // @[Cat.scala 29:58]
  assign _T_516 = _T_511 ? _T_515 : _T_503; // @[Shift.scala 91:22]
  assign _T_517 = _T_506[2:0]; // @[Shift.scala 92:77]
  assign _T_518 = _T_516[14:4]; // @[Shift.scala 90:30]
  assign _T_519 = _T_516[3:0]; // @[Shift.scala 90:48]
  assign _T_520 = _T_519 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{10'd0}, _T_520}; // @[Shift.scala 90:39]
  assign _T_521 = _T_518 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_522 = _T_517[2]; // @[Shift.scala 12:21]
  assign _T_523 = _T_516[14]; // @[Shift.scala 12:21]
  assign _T_525 = _T_523 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_526 = {_T_525,_T_521}; // @[Cat.scala 29:58]
  assign _T_527 = _T_522 ? _T_526 : _T_516; // @[Shift.scala 91:22]
  assign _T_528 = _T_517[1:0]; // @[Shift.scala 92:77]
  assign _T_529 = _T_527[14:2]; // @[Shift.scala 90:30]
  assign _T_530 = _T_527[1:0]; // @[Shift.scala 90:48]
  assign _T_531 = _T_530 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_8 = {{12'd0}, _T_531}; // @[Shift.scala 90:39]
  assign _T_532 = _T_529 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_533 = _T_528[1]; // @[Shift.scala 12:21]
  assign _T_534 = _T_527[14]; // @[Shift.scala 12:21]
  assign _T_536 = _T_534 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_537 = {_T_536,_T_532}; // @[Cat.scala 29:58]
  assign _T_538 = _T_533 ? _T_537 : _T_527; // @[Shift.scala 91:22]
  assign _T_539 = _T_528[0:0]; // @[Shift.scala 92:77]
  assign _T_540 = _T_538[14:1]; // @[Shift.scala 90:30]
  assign _T_541 = _T_538[0:0]; // @[Shift.scala 90:48]
  assign _GEN_9 = {{13'd0}, _T_541}; // @[Shift.scala 90:39]
  assign _T_543 = _T_540 | _GEN_9; // @[Shift.scala 90:39]
  assign _T_545 = _T_538[14]; // @[Shift.scala 12:21]
  assign _T_546 = {_T_545,_T_543}; // @[Cat.scala 29:58]
  assign _T_547 = _T_539 ? _T_546 : _T_538; // @[Shift.scala 91:22]
  assign _T_550 = _T_512 ? 15'h7fff : 15'h0; // @[Bitwise.scala 71:12]
  assign _T_551 = _T_505 ? _T_547 : _T_550; // @[Shift.scala 39:10]
  assign _T_552 = _T_551[3]; // @[convert.scala 55:31]
  assign _T_553 = _T_551[2]; // @[convert.scala 56:31]
  assign _T_554 = _T_551[1]; // @[convert.scala 57:31]
  assign _T_555 = _T_551[0]; // @[convert.scala 58:31]
  assign _T_556 = _T_551[14:3]; // @[convert.scala 59:69]
  assign _T_557 = _T_556 != 12'h0; // @[convert.scala 59:81]
  assign _T_558 = ~ _T_557; // @[convert.scala 59:50]
  assign _T_560 = _T_556 == 12'hfff; // @[convert.scala 60:81]
  assign _T_561 = _T_552 | _T_554; // @[convert.scala 61:44]
  assign _T_562 = _T_561 | _T_555; // @[convert.scala 61:52]
  assign _T_563 = _T_553 & _T_562; // @[convert.scala 61:36]
  assign _T_564 = ~ _T_560; // @[convert.scala 62:63]
  assign _T_565 = _T_564 & _T_563; // @[convert.scala 62:103]
  assign _T_566 = _T_558 | _T_565; // @[convert.scala 62:60]
  assign _GEN_10 = {{11'd0}, _T_566}; // @[convert.scala 63:56]
  assign _T_569 = _T_556 + _GEN_10; // @[convert.scala 63:56]
  assign _T_570 = {sumSign,_T_569}; // @[Cat.scala 29:58]
  assign _T_572 = decS_isZero ? 13'h0 : _T_570; // @[Mux.scala 87:16]
  assign io_S = decS_isNaR ? 13'h1000 : _T_572; // @[PositAdder.scala 56:8]
endmodule
