module PositDivSqrter8_2(
  input        clock,
  input        reset,
  output       io_inReady,
  input        io_inValid,
  input        io_sqrtOp,
  input  [7:0] io_A,
  input  [7:0] io_B,
  output       io_diviValid,
  output       io_sqrtValid,
  output       io_invalidExc,
  output [7:0] io_Q
);
  reg [2:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [6:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [2:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [6:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [6:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [5:0] _T_4; // @[convert.scala 19:24]
  wire [5:0] _T_5; // @[convert.scala 19:43]
  wire [5:0] _T_6; // @[convert.scala 19:39]
  wire [3:0] _T_7; // @[LZD.scala 43:32]
  wire [1:0] _T_8; // @[LZD.scala 43:32]
  wire  _T_9; // @[LZD.scala 39:14]
  wire  _T_10; // @[LZD.scala 39:21]
  wire  _T_11; // @[LZD.scala 39:30]
  wire  _T_12; // @[LZD.scala 39:27]
  wire  _T_13; // @[LZD.scala 39:25]
  wire [1:0] _T_14; // @[Cat.scala 29:58]
  wire [1:0] _T_15; // @[LZD.scala 44:32]
  wire  _T_16; // @[LZD.scala 39:14]
  wire  _T_17; // @[LZD.scala 39:21]
  wire  _T_18; // @[LZD.scala 39:30]
  wire  _T_19; // @[LZD.scala 39:27]
  wire  _T_20; // @[LZD.scala 39:25]
  wire [1:0] _T_21; // @[Cat.scala 29:58]
  wire  _T_22; // @[Shift.scala 12:21]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[LZD.scala 49:16]
  wire  _T_25; // @[LZD.scala 49:27]
  wire  _T_26; // @[LZD.scala 49:25]
  wire  _T_27; // @[LZD.scala 49:47]
  wire  _T_28; // @[LZD.scala 49:59]
  wire  _T_29; // @[LZD.scala 49:35]
  wire [2:0] _T_31; // @[Cat.scala 29:58]
  wire [1:0] _T_32; // @[LZD.scala 44:32]
  wire  _T_33; // @[LZD.scala 39:14]
  wire  _T_34; // @[LZD.scala 39:21]
  wire  _T_35; // @[LZD.scala 39:30]
  wire  _T_36; // @[LZD.scala 39:27]
  wire  _T_37; // @[LZD.scala 39:25]
  wire [1:0] _T_38; // @[Cat.scala 29:58]
  wire  _T_39; // @[Shift.scala 12:21]
  wire [1:0] _T_41; // @[LZD.scala 55:32]
  wire [1:0] _T_42; // @[LZD.scala 55:20]
  wire [2:0] _T_43; // @[Cat.scala 29:58]
  wire [2:0] _T_44; // @[convert.scala 21:22]
  wire [4:0] _T_45; // @[convert.scala 22:36]
  wire  _T_46; // @[Shift.scala 16:24]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 64:52]
  wire [4:0] _T_51; // @[Cat.scala 29:58]
  wire [4:0] _T_52; // @[Shift.scala 64:27]
  wire [1:0] _T_53; // @[Shift.scala 66:70]
  wire  _T_54; // @[Shift.scala 12:21]
  wire [2:0] _T_55; // @[Shift.scala 64:52]
  wire [4:0] _T_57; // @[Cat.scala 29:58]
  wire [4:0] _T_58; // @[Shift.scala 64:27]
  wire  _T_59; // @[Shift.scala 66:70]
  wire [3:0] _T_61; // @[Shift.scala 64:52]
  wire [4:0] _T_62; // @[Cat.scala 29:58]
  wire [4:0] _T_63; // @[Shift.scala 64:27]
  wire [4:0] _T_64; // @[Shift.scala 16:10]
  wire [1:0] _T_65; // @[convert.scala 23:34]
  wire [2:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_67; // @[convert.scala 25:26]
  wire [2:0] _T_69; // @[convert.scala 25:42]
  wire [1:0] _T_72; // @[convert.scala 26:67]
  wire [1:0] _T_73; // @[convert.scala 26:51]
  wire [5:0] _T_74; // @[Cat.scala 29:58]
  wire [6:0] _T_76; // @[convert.scala 29:56]
  wire  _T_77; // @[convert.scala 29:60]
  wire  _T_78; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_81; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_90; // @[convert.scala 18:24]
  wire  _T_91; // @[convert.scala 18:40]
  wire  _T_92; // @[convert.scala 18:36]
  wire [5:0] _T_93; // @[convert.scala 19:24]
  wire [5:0] _T_94; // @[convert.scala 19:43]
  wire [5:0] _T_95; // @[convert.scala 19:39]
  wire [3:0] _T_96; // @[LZD.scala 43:32]
  wire [1:0] _T_97; // @[LZD.scala 43:32]
  wire  _T_98; // @[LZD.scala 39:14]
  wire  _T_99; // @[LZD.scala 39:21]
  wire  _T_100; // @[LZD.scala 39:30]
  wire  _T_101; // @[LZD.scala 39:27]
  wire  _T_102; // @[LZD.scala 39:25]
  wire [1:0] _T_103; // @[Cat.scala 29:58]
  wire [1:0] _T_104; // @[LZD.scala 44:32]
  wire  _T_105; // @[LZD.scala 39:14]
  wire  _T_106; // @[LZD.scala 39:21]
  wire  _T_107; // @[LZD.scala 39:30]
  wire  _T_108; // @[LZD.scala 39:27]
  wire  _T_109; // @[LZD.scala 39:25]
  wire [1:0] _T_110; // @[Cat.scala 29:58]
  wire  _T_111; // @[Shift.scala 12:21]
  wire  _T_112; // @[Shift.scala 12:21]
  wire  _T_113; // @[LZD.scala 49:16]
  wire  _T_114; // @[LZD.scala 49:27]
  wire  _T_115; // @[LZD.scala 49:25]
  wire  _T_116; // @[LZD.scala 49:47]
  wire  _T_117; // @[LZD.scala 49:59]
  wire  _T_118; // @[LZD.scala 49:35]
  wire [2:0] _T_120; // @[Cat.scala 29:58]
  wire [1:0] _T_121; // @[LZD.scala 44:32]
  wire  _T_122; // @[LZD.scala 39:14]
  wire  _T_123; // @[LZD.scala 39:21]
  wire  _T_124; // @[LZD.scala 39:30]
  wire  _T_125; // @[LZD.scala 39:27]
  wire  _T_126; // @[LZD.scala 39:25]
  wire [1:0] _T_127; // @[Cat.scala 29:58]
  wire  _T_128; // @[Shift.scala 12:21]
  wire [1:0] _T_130; // @[LZD.scala 55:32]
  wire [1:0] _T_131; // @[LZD.scala 55:20]
  wire [2:0] _T_132; // @[Cat.scala 29:58]
  wire [2:0] _T_133; // @[convert.scala 21:22]
  wire [4:0] _T_134; // @[convert.scala 22:36]
  wire  _T_135; // @[Shift.scala 16:24]
  wire  _T_137; // @[Shift.scala 12:21]
  wire  _T_138; // @[Shift.scala 64:52]
  wire [4:0] _T_140; // @[Cat.scala 29:58]
  wire [4:0] _T_141; // @[Shift.scala 64:27]
  wire [1:0] _T_142; // @[Shift.scala 66:70]
  wire  _T_143; // @[Shift.scala 12:21]
  wire [2:0] _T_144; // @[Shift.scala 64:52]
  wire [4:0] _T_146; // @[Cat.scala 29:58]
  wire [4:0] _T_147; // @[Shift.scala 64:27]
  wire  _T_148; // @[Shift.scala 66:70]
  wire [3:0] _T_150; // @[Shift.scala 64:52]
  wire [4:0] _T_151; // @[Cat.scala 29:58]
  wire [4:0] _T_152; // @[Shift.scala 64:27]
  wire [4:0] _T_153; // @[Shift.scala 16:10]
  wire [1:0] _T_154; // @[convert.scala 23:34]
  wire [2:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_156; // @[convert.scala 25:26]
  wire [2:0] _T_158; // @[convert.scala 25:42]
  wire [1:0] _T_161; // @[convert.scala 26:67]
  wire [1:0] _T_162; // @[convert.scala 26:51]
  wire [5:0] _T_163; // @[Cat.scala 29:58]
  wire [6:0] _T_165; // @[convert.scala 29:56]
  wire  _T_166; // @[convert.scala 29:60]
  wire  _T_167; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_170; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_179; // @[Bitwise.scala 71:12]
  wire  _T_180; // @[PositDivisionSqrt.scala 80:40]
  wire [6:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_182; // @[PositDivisionSqrt.scala 82:31]
  wire [6:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_185; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_186; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_187; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_188; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_189; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_190; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_191; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_192; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_193; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_194; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [6:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_197; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_198; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_199; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_200; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_201; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_202; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_203; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_204; // @[PositDivisionSqrt.scala 117:30]
  wire [2:0] _T_206; // @[PositDivisionSqrt.scala 119:26]
  wire [2:0] _T_207; // @[PositDivisionSqrt.scala 118:20]
  wire [2:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [2:0] _T_208; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_210; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_211; // @[PositDivisionSqrt.scala 123:27]
  wire [2:0] _T_213; // @[PositDivisionSqrt.scala 123:52]
  wire [2:0] _T_214; // @[PositDivisionSqrt.scala 123:20]
  wire [2:0] _T_215; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_217; // @[PositDivisionSqrt.scala 124:27]
  wire [2:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [2:0] _T_219; // @[PositDivisionSqrt.scala 123:64]
  wire [4:0] _T_220; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_222; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_223; // @[PositDivisionSqrt.scala 137:28]
  wire [7:0] _T_224; // @[PositDivisionSqrt.scala 146:22]
  wire [5:0] bitMask; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_226; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_227; // @[PositDivisionSqrt.scala 148:23]
  wire [6:0] _T_228; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_229; // @[PositDivisionSqrt.scala 149:23]
  wire [7:0] _T_230; // @[PositDivisionSqrt.scala 149:46]
  wire [6:0] _T_231; // @[PositDivisionSqrt.scala 149:56]
  wire [6:0] _T_232; // @[PositDivisionSqrt.scala 149:16]
  wire [6:0] _T_233; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_234; // @[PositDivisionSqrt.scala 150:17]
  wire [6:0] _T_235; // @[PositDivisionSqrt.scala 150:16]
  wire [6:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_237; // @[PositDivisionSqrt.scala 152:29]
  wire [6:0] _T_238; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_239; // @[PositDivisionSqrt.scala 153:29]
  wire [3:0] _T_240; // @[PositDivisionSqrt.scala 153:22]
  wire [6:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [6:0] _T_241; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_243; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_244; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_245; // @[PositDivisionSqrt.scala 154:57]
  wire [6:0] _T_248; // @[Cat.scala 29:58]
  wire [6:0] _T_249; // @[PositDivisionSqrt.scala 154:22]
  wire [6:0] _T_250; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_252; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_253; // @[PositDivisionSqrt.scala 156:79]
  wire [2:0] _T_255; // @[Bitwise.scala 71:12]
  wire [5:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [5:0] _T_256; // @[PositDivisionSqrt.scala 156:53]
  wire [6:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [6:0] _T_257; // @[PositDivisionSqrt.scala 155:51]
  wire [4:0] _T_258; // @[PositDivisionSqrt.scala 157:53]
  wire [6:0] _GEN_14; // @[PositDivisionSqrt.scala 156:85]
  wire [6:0] _T_259; // @[PositDivisionSqrt.scala 156:85]
  wire [6:0] _T_260; // @[PositDivisionSqrt.scala 155:22]
  wire [6:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_262; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_263; // @[PositDivisionSqrt.scala 162:40]
  wire [6:0] _T_266; // @[PositDivisionSqrt.scala 163:97]
  wire [6:0] _T_268; // @[PositDivisionSqrt.scala 164:97]
  wire [6:0] _T_269; // @[PositDivisionSqrt.scala 161:92]
  wire [7:0] _T_274; // @[PositDivisionSqrt.scala 168:98]
  wire [6:0] _T_275; // @[PositDivisionSqrt.scala 168:108]
  wire [6:0] _T_277; // @[PositDivisionSqrt.scala 168:112]
  wire [6:0] _T_281; // @[PositDivisionSqrt.scala 169:112]
  wire [6:0] _T_282; // @[PositDivisionSqrt.scala 166:26]
  wire [6:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_283; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_284; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_286; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_287; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_288; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_289; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_290; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_292; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_293; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_294; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_295; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_296; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_299; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_300; // @[PositDivisionSqrt.scala 187:28]
  wire [6:0] _T_303; // @[PositDivisionSqrt.scala 188:47]
  wire [6:0] _T_304; // @[PositDivisionSqrt.scala 188:18]
  wire [4:0] _T_306; // @[PositDivisionSqrt.scala 189:18]
  wire [6:0] _GEN_15; // @[PositDivisionSqrt.scala 188:72]
  wire [6:0] _T_307; // @[PositDivisionSqrt.scala 188:72]
  wire [6:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [6:0] _T_309; // @[PositDivisionSqrt.scala 190:47]
  wire [6:0] _T_310; // @[PositDivisionSqrt.scala 190:18]
  wire [6:0] _T_311; // @[PositDivisionSqrt.scala 189:72]
  wire [1:0] _T_313; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [6:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [6:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [2:0] _T_316; // @[PositDivisionSqrt.scala 200:97]
  wire [2:0] _T_317; // @[PositDivisionSqrt.scala 201:97]
  wire [2:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_318; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_319; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_320; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_322; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_323; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_324; // @[Cat.scala 29:58]
  wire [2:0] _T_325; // @[PositDivisionSqrt.scala 209:63]
  wire [6:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] _T_327; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [6:0] _T_329; // @[Mux.scala 87:16]
  wire [6:0] _T_330; // @[Mux.scala 87:16]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [5:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [5:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [1:0] _T_335; // @[convert.scala 46:61]
  wire [1:0] _T_336; // @[convert.scala 46:52]
  wire [1:0] _T_338; // @[convert.scala 46:42]
  wire [3:0] _T_339; // @[convert.scala 48:34]
  wire  _T_340; // @[convert.scala 49:36]
  wire [3:0] _T_342; // @[convert.scala 50:36]
  wire [3:0] _T_343; // @[convert.scala 50:36]
  wire [3:0] _T_344; // @[convert.scala 50:28]
  wire  _T_345; // @[convert.scala 51:31]
  wire  _T_346; // @[convert.scala 52:43]
  wire [9:0] _T_350; // @[Cat.scala 29:58]
  wire [3:0] _T_351; // @[Shift.scala 39:17]
  wire  _T_352; // @[Shift.scala 39:24]
  wire [1:0] _T_354; // @[Shift.scala 90:30]
  wire [7:0] _T_355; // @[Shift.scala 90:48]
  wire  _T_356; // @[Shift.scala 90:57]
  wire [1:0] _GEN_20; // @[Shift.scala 90:39]
  wire [1:0] _T_357; // @[Shift.scala 90:39]
  wire  _T_358; // @[Shift.scala 12:21]
  wire  _T_359; // @[Shift.scala 12:21]
  wire [7:0] _T_361; // @[Bitwise.scala 71:12]
  wire [9:0] _T_362; // @[Cat.scala 29:58]
  wire [9:0] _T_363; // @[Shift.scala 91:22]
  wire [2:0] _T_364; // @[Shift.scala 92:77]
  wire [5:0] _T_365; // @[Shift.scala 90:30]
  wire [3:0] _T_366; // @[Shift.scala 90:48]
  wire  _T_367; // @[Shift.scala 90:57]
  wire [5:0] _GEN_21; // @[Shift.scala 90:39]
  wire [5:0] _T_368; // @[Shift.scala 90:39]
  wire  _T_369; // @[Shift.scala 12:21]
  wire  _T_370; // @[Shift.scala 12:21]
  wire [3:0] _T_372; // @[Bitwise.scala 71:12]
  wire [9:0] _T_373; // @[Cat.scala 29:58]
  wire [9:0] _T_374; // @[Shift.scala 91:22]
  wire [1:0] _T_375; // @[Shift.scala 92:77]
  wire [7:0] _T_376; // @[Shift.scala 90:30]
  wire [1:0] _T_377; // @[Shift.scala 90:48]
  wire  _T_378; // @[Shift.scala 90:57]
  wire [7:0] _GEN_22; // @[Shift.scala 90:39]
  wire [7:0] _T_379; // @[Shift.scala 90:39]
  wire  _T_380; // @[Shift.scala 12:21]
  wire  _T_381; // @[Shift.scala 12:21]
  wire [1:0] _T_383; // @[Bitwise.scala 71:12]
  wire [9:0] _T_384; // @[Cat.scala 29:58]
  wire [9:0] _T_385; // @[Shift.scala 91:22]
  wire  _T_386; // @[Shift.scala 92:77]
  wire [8:0] _T_387; // @[Shift.scala 90:30]
  wire  _T_388; // @[Shift.scala 90:48]
  wire [8:0] _GEN_23; // @[Shift.scala 90:39]
  wire [8:0] _T_390; // @[Shift.scala 90:39]
  wire  _T_392; // @[Shift.scala 12:21]
  wire [9:0] _T_393; // @[Cat.scala 29:58]
  wire [9:0] _T_394; // @[Shift.scala 91:22]
  wire [9:0] _T_397; // @[Bitwise.scala 71:12]
  wire [9:0] _T_398; // @[Shift.scala 39:10]
  wire  _T_399; // @[convert.scala 55:31]
  wire  _T_400; // @[convert.scala 56:31]
  wire  _T_401; // @[convert.scala 57:31]
  wire  _T_402; // @[convert.scala 58:31]
  wire [6:0] _T_403; // @[convert.scala 59:69]
  wire  _T_404; // @[convert.scala 59:81]
  wire  _T_405; // @[convert.scala 59:50]
  wire  _T_407; // @[convert.scala 60:81]
  wire  _T_408; // @[convert.scala 61:44]
  wire  _T_409; // @[convert.scala 61:52]
  wire  _T_410; // @[convert.scala 61:36]
  wire  _T_411; // @[convert.scala 62:63]
  wire  _T_412; // @[convert.scala 62:103]
  wire  _T_413; // @[convert.scala 62:60]
  wire [6:0] _GEN_24; // @[convert.scala 63:56]
  wire [6:0] _T_416; // @[convert.scala 63:56]
  wire [7:0] _T_417; // @[Cat.scala 29:58]
  wire [7:0] _T_419; // @[Mux.scala 87:16]
  assign _T_1 = io_A[7]; // @[convert.scala 18:24]
  assign _T_2 = io_A[6]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[6:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[5:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[5:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[3:2]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8 != 2'h0; // @[LZD.scala 39:14]
  assign _T_10 = _T_8[1]; // @[LZD.scala 39:21]
  assign _T_11 = _T_8[0]; // @[LZD.scala 39:30]
  assign _T_12 = ~ _T_11; // @[LZD.scala 39:27]
  assign _T_13 = _T_10 | _T_12; // @[LZD.scala 39:25]
  assign _T_14 = {_T_9,_T_13}; // @[Cat.scala 29:58]
  assign _T_15 = _T_7[1:0]; // @[LZD.scala 44:32]
  assign _T_16 = _T_15 != 2'h0; // @[LZD.scala 39:14]
  assign _T_17 = _T_15[1]; // @[LZD.scala 39:21]
  assign _T_18 = _T_15[0]; // @[LZD.scala 39:30]
  assign _T_19 = ~ _T_18; // @[LZD.scala 39:27]
  assign _T_20 = _T_17 | _T_19; // @[LZD.scala 39:25]
  assign _T_21 = {_T_16,_T_20}; // @[Cat.scala 29:58]
  assign _T_22 = _T_14[1]; // @[Shift.scala 12:21]
  assign _T_23 = _T_21[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22 | _T_23; // @[LZD.scala 49:16]
  assign _T_25 = ~ _T_23; // @[LZD.scala 49:27]
  assign _T_26 = _T_22 | _T_25; // @[LZD.scala 49:25]
  assign _T_27 = _T_14[0:0]; // @[LZD.scala 49:47]
  assign _T_28 = _T_21[0:0]; // @[LZD.scala 49:59]
  assign _T_29 = _T_22 ? _T_27 : _T_28; // @[LZD.scala 49:35]
  assign _T_31 = {_T_24,_T_26,_T_29}; // @[Cat.scala 29:58]
  assign _T_32 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_33 = _T_32 != 2'h0; // @[LZD.scala 39:14]
  assign _T_34 = _T_32[1]; // @[LZD.scala 39:21]
  assign _T_35 = _T_32[0]; // @[LZD.scala 39:30]
  assign _T_36 = ~ _T_35; // @[LZD.scala 39:27]
  assign _T_37 = _T_34 | _T_36; // @[LZD.scala 39:25]
  assign _T_38 = {_T_33,_T_37}; // @[Cat.scala 29:58]
  assign _T_39 = _T_31[2]; // @[Shift.scala 12:21]
  assign _T_41 = _T_31[1:0]; // @[LZD.scala 55:32]
  assign _T_42 = _T_39 ? _T_41 : _T_38; // @[LZD.scala 55:20]
  assign _T_43 = {_T_39,_T_42}; // @[Cat.scala 29:58]
  assign _T_44 = ~ _T_43; // @[convert.scala 21:22]
  assign _T_45 = io_A[4:0]; // @[convert.scala 22:36]
  assign _T_46 = _T_44 < 3'h5; // @[Shift.scala 16:24]
  assign _T_48 = _T_44[2]; // @[Shift.scala 12:21]
  assign _T_49 = _T_45[0:0]; // @[Shift.scala 64:52]
  assign _T_51 = {_T_49,4'h0}; // @[Cat.scala 29:58]
  assign _T_52 = _T_48 ? _T_51 : _T_45; // @[Shift.scala 64:27]
  assign _T_53 = _T_44[1:0]; // @[Shift.scala 66:70]
  assign _T_54 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_55 = _T_52[2:0]; // @[Shift.scala 64:52]
  assign _T_57 = {_T_55,2'h0}; // @[Cat.scala 29:58]
  assign _T_58 = _T_54 ? _T_57 : _T_52; // @[Shift.scala 64:27]
  assign _T_59 = _T_53[0:0]; // @[Shift.scala 66:70]
  assign _T_61 = _T_58[3:0]; // @[Shift.scala 64:52]
  assign _T_62 = {_T_61,1'h0}; // @[Cat.scala 29:58]
  assign _T_63 = _T_59 ? _T_62 : _T_58; // @[Shift.scala 64:27]
  assign _T_64 = _T_46 ? _T_63 : 5'h0; // @[Shift.scala 16:10]
  assign _T_65 = _T_64[4:3]; // @[convert.scala 23:34]
  assign decA_fraction = _T_64[2:0]; // @[convert.scala 24:34]
  assign _T_67 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_69 = _T_3 ? _T_44 : _T_43; // @[convert.scala 25:42]
  assign _T_72 = ~ _T_65; // @[convert.scala 26:67]
  assign _T_73 = _T_1 ? _T_72 : _T_65; // @[convert.scala 26:51]
  assign _T_74 = {_T_67,_T_69,_T_73}; // @[Cat.scala 29:58]
  assign _T_76 = io_A[6:0]; // @[convert.scala 29:56]
  assign _T_77 = _T_76 != 7'h0; // @[convert.scala 29:60]
  assign _T_78 = ~ _T_77; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_78; // @[convert.scala 29:39]
  assign _T_81 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_81 & _T_78; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_74); // @[convert.scala 32:24]
  assign _T_90 = io_B[7]; // @[convert.scala 18:24]
  assign _T_91 = io_B[6]; // @[convert.scala 18:40]
  assign _T_92 = _T_90 ^ _T_91; // @[convert.scala 18:36]
  assign _T_93 = io_B[6:1]; // @[convert.scala 19:24]
  assign _T_94 = io_B[5:0]; // @[convert.scala 19:43]
  assign _T_95 = _T_93 ^ _T_94; // @[convert.scala 19:39]
  assign _T_96 = _T_95[5:2]; // @[LZD.scala 43:32]
  assign _T_97 = _T_96[3:2]; // @[LZD.scala 43:32]
  assign _T_98 = _T_97 != 2'h0; // @[LZD.scala 39:14]
  assign _T_99 = _T_97[1]; // @[LZD.scala 39:21]
  assign _T_100 = _T_97[0]; // @[LZD.scala 39:30]
  assign _T_101 = ~ _T_100; // @[LZD.scala 39:27]
  assign _T_102 = _T_99 | _T_101; // @[LZD.scala 39:25]
  assign _T_103 = {_T_98,_T_102}; // @[Cat.scala 29:58]
  assign _T_104 = _T_96[1:0]; // @[LZD.scala 44:32]
  assign _T_105 = _T_104 != 2'h0; // @[LZD.scala 39:14]
  assign _T_106 = _T_104[1]; // @[LZD.scala 39:21]
  assign _T_107 = _T_104[0]; // @[LZD.scala 39:30]
  assign _T_108 = ~ _T_107; // @[LZD.scala 39:27]
  assign _T_109 = _T_106 | _T_108; // @[LZD.scala 39:25]
  assign _T_110 = {_T_105,_T_109}; // @[Cat.scala 29:58]
  assign _T_111 = _T_103[1]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110[1]; // @[Shift.scala 12:21]
  assign _T_113 = _T_111 | _T_112; // @[LZD.scala 49:16]
  assign _T_114 = ~ _T_112; // @[LZD.scala 49:27]
  assign _T_115 = _T_111 | _T_114; // @[LZD.scala 49:25]
  assign _T_116 = _T_103[0:0]; // @[LZD.scala 49:47]
  assign _T_117 = _T_110[0:0]; // @[LZD.scala 49:59]
  assign _T_118 = _T_111 ? _T_116 : _T_117; // @[LZD.scala 49:35]
  assign _T_120 = {_T_113,_T_115,_T_118}; // @[Cat.scala 29:58]
  assign _T_121 = _T_95[1:0]; // @[LZD.scala 44:32]
  assign _T_122 = _T_121 != 2'h0; // @[LZD.scala 39:14]
  assign _T_123 = _T_121[1]; // @[LZD.scala 39:21]
  assign _T_124 = _T_121[0]; // @[LZD.scala 39:30]
  assign _T_125 = ~ _T_124; // @[LZD.scala 39:27]
  assign _T_126 = _T_123 | _T_125; // @[LZD.scala 39:25]
  assign _T_127 = {_T_122,_T_126}; // @[Cat.scala 29:58]
  assign _T_128 = _T_120[2]; // @[Shift.scala 12:21]
  assign _T_130 = _T_120[1:0]; // @[LZD.scala 55:32]
  assign _T_131 = _T_128 ? _T_130 : _T_127; // @[LZD.scala 55:20]
  assign _T_132 = {_T_128,_T_131}; // @[Cat.scala 29:58]
  assign _T_133 = ~ _T_132; // @[convert.scala 21:22]
  assign _T_134 = io_B[4:0]; // @[convert.scala 22:36]
  assign _T_135 = _T_133 < 3'h5; // @[Shift.scala 16:24]
  assign _T_137 = _T_133[2]; // @[Shift.scala 12:21]
  assign _T_138 = _T_134[0:0]; // @[Shift.scala 64:52]
  assign _T_140 = {_T_138,4'h0}; // @[Cat.scala 29:58]
  assign _T_141 = _T_137 ? _T_140 : _T_134; // @[Shift.scala 64:27]
  assign _T_142 = _T_133[1:0]; // @[Shift.scala 66:70]
  assign _T_143 = _T_142[1]; // @[Shift.scala 12:21]
  assign _T_144 = _T_141[2:0]; // @[Shift.scala 64:52]
  assign _T_146 = {_T_144,2'h0}; // @[Cat.scala 29:58]
  assign _T_147 = _T_143 ? _T_146 : _T_141; // @[Shift.scala 64:27]
  assign _T_148 = _T_142[0:0]; // @[Shift.scala 66:70]
  assign _T_150 = _T_147[3:0]; // @[Shift.scala 64:52]
  assign _T_151 = {_T_150,1'h0}; // @[Cat.scala 29:58]
  assign _T_152 = _T_148 ? _T_151 : _T_147; // @[Shift.scala 64:27]
  assign _T_153 = _T_135 ? _T_152 : 5'h0; // @[Shift.scala 16:10]
  assign _T_154 = _T_153[4:3]; // @[convert.scala 23:34]
  assign decB_fraction = _T_153[2:0]; // @[convert.scala 24:34]
  assign _T_156 = _T_92 == 1'h0; // @[convert.scala 25:26]
  assign _T_158 = _T_92 ? _T_133 : _T_132; // @[convert.scala 25:42]
  assign _T_161 = ~ _T_154; // @[convert.scala 26:67]
  assign _T_162 = _T_90 ? _T_161 : _T_154; // @[convert.scala 26:51]
  assign _T_163 = {_T_156,_T_158,_T_162}; // @[Cat.scala 29:58]
  assign _T_165 = io_B[6:0]; // @[convert.scala 29:56]
  assign _T_166 = _T_165 != 7'h0; // @[convert.scala 29:60]
  assign _T_167 = ~ _T_166; // @[convert.scala 29:41]
  assign decB_isNaR = _T_90 & _T_167; // @[convert.scala 29:39]
  assign _T_170 = _T_90 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_170 & _T_167; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_163); // @[convert.scala 32:24]
  assign _T_179 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_180 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_179,_T_180,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_182 = ~ _T_90; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_90,_T_182,decB_fraction,2'h0}; // @[Cat.scala 29:58]
  assign _T_185 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_185 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_186 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_187 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_188 = _T_187 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_189 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_190 = decA_isZero & _T_189; // @[PositDivisionSqrt.scala 94:43]
  assign _T_191 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_192 = _T_190 & _T_191; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_193 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_194 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_193 & _T_194; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_193 & _T_81; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_197 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_197; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 3'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 3'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_198 = sigX_Z[6]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_199 = sigX_Z[4]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_198 ^ _T_199; // @[PositDivisionSqrt.scala 113:50]
  assign _T_200 = cycleNum == 3'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_200 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_201 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_202 = _T_201 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_203 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_204 = entering & _T_203; // @[PositDivisionSqrt.scala 117:30]
  assign _T_206 = io_sqrtOp ? 3'h5 : 3'h7; // @[PositDivisionSqrt.scala 119:26]
  assign _T_207 = entering_normalCase ? _T_206 : 3'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{2'd0}, _T_204}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_208 = _GEN_9 | _T_207; // @[PositDivisionSqrt.scala 117:64]
  assign _T_210 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_211 = _T_201 & _T_210; // @[PositDivisionSqrt.scala 123:27]
  assign _T_213 = cycleNum - 3'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_214 = _T_211 ? _T_213 : 3'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_215 = _T_208 | _T_214; // @[PositDivisionSqrt.scala 122:64]
  assign _T_217 = _T_201 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{2'd0}, _T_217}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_219 = _T_215 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_220 = decA_scale[5:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_222 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_223 = entering_normalCase & _T_222; // @[PositDivisionSqrt.scala 137:28]
  assign _T_224 = 8'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign bitMask = _T_224[7:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_226 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_227 = ready & _T_226; // @[PositDivisionSqrt.scala 148:23]
  assign _T_228 = _T_227 ? sigA_S : 7'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_229 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_230 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_231 = _T_230[6:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_232 = _T_229 ? _T_231 : 7'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_233 = _T_228 | _T_232; // @[PositDivisionSqrt.scala 148:66]
  assign _T_234 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_235 = _T_234 ? rem_Z : 7'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_233 | _T_235; // @[PositDivisionSqrt.scala 149:66]
  assign _T_237 = ready & _T_222; // @[PositDivisionSqrt.scala 152:29]
  assign _T_238 = _T_237 ? sigB_S : 7'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_239 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_240 = _T_239 ? 4'h8 : 4'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_240}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_241 = _T_238 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_243 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_244 = _T_234 & _T_243; // @[PositDivisionSqrt.scala 154:30]
  assign _T_245 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_248 = {signB_Z,_T_245,fractB_Z,2'h0}; // @[Cat.scala 29:58]
  assign _T_249 = _T_244 ? _T_248 : 7'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_250 = _T_241 | _T_249; // @[PositDivisionSqrt.scala 153:93]
  assign _T_252 = _T_234 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_253 = rem[6:6]; // @[PositDivisionSqrt.scala 156:79]
  assign _T_255 = _T_253 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _GEN_12 = {{3'd0}, _T_255}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_256 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_256}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_257 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_258 = bitMask[5:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_258}; // @[PositDivisionSqrt.scala 156:85]
  assign _T_259 = _T_257 | _GEN_14; // @[PositDivisionSqrt.scala 156:85]
  assign _T_260 = _T_252 ? _T_259 : 7'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_250 | _T_260; // @[PositDivisionSqrt.scala 154:93]
  assign _T_262 = trialTerm[6:6]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_263 = _T_253 ^ _T_262; // @[PositDivisionSqrt.scala 162:40]
  assign _T_266 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_268 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_269 = _T_263 ? _T_266 : _T_268; // @[PositDivisionSqrt.scala 161:92]
  assign _T_274 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_275 = _T_274[6:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_277 = _T_275 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_281 = _T_275 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_282 = _T_263 ? _T_277 : _T_281; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_269 : _T_282; // @[PositDivisionSqrt.scala 159:27]
  assign _T_283 = trialRem != 7'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_283 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_284 = rem != 7'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_284 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_286 = trialRem[6:6]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_287 = _T_262 ^ _T_286; // @[PositDivisionSqrt.scala 176:49]
  assign _T_288 = ~ _T_287; // @[PositDivisionSqrt.scala 176:29]
  assign _T_289 = sigX_Z[6:6]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_290 = ~ _T_289; // @[PositDivisionSqrt.scala 178:49]
  assign _T_292 = remIsZero ? _T_289 : _T_288; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_290 : _T_292; // @[Mux.scala 87:16]
  assign _T_293 = cycleNum > 3'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_294 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_295 = _T_293 & _T_294; // @[PositDivisionSqrt.scala 183:48]
  assign _T_296 = entering_normalCase | _T_295; // @[PositDivisionSqrt.scala 183:28]
  assign _T_299 = _T_234 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_300 = entering_normalCase | _T_299; // @[PositDivisionSqrt.scala 187:28]
  assign _T_303 = {newBit, 6'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_304 = _T_237 ? _T_303 : 7'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_306 = _T_239 ? 5'h10 : 5'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_306}; // @[PositDivisionSqrt.scala 188:72]
  assign _T_307 = _T_304 | _GEN_15; // @[PositDivisionSqrt.scala 188:72]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_309 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_310 = _T_234 ? _T_309 : 7'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_311 = _T_307 | _T_310; // @[PositDivisionSqrt.scala 189:72]
  assign _T_313 = {_T_289, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_313 : {{1'd0}, _T_289}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{5'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_316 = realSigX[3:1]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_317 = realSigX[2:0]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_316 : _T_317; // @[PositDivisionSqrt.scala 198:21]
  assign _T_318 = realSigX[6]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_319 = realSigX[4]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_320 = _T_318 ^ _T_319; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_320; // @[PositDivisionSqrt.scala 205:23]
  assign _T_322 = realSigX[3]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_318 ^ _T_322; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_323 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_323; // @[PositDivisionSqrt.scala 208:36]
  assign _T_324 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_325 = {1'b0,$signed(_T_324)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{4{_T_325[2]}},_T_325}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_327 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_327); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-7'sh18); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(7'sh18); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[6:6]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_329 = underflow ? $signed(-7'sh18) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_330 = overflow ? $signed(7'sh18) : $signed(_T_329); // @[Mux.scala 87:16]
  assign outValid = cycleNum == 3'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_330[5:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_335 = decQ_scale[1:0]; // @[convert.scala 46:61]
  assign _T_336 = ~ _T_335; // @[convert.scala 46:52]
  assign _T_338 = decQ_sign ? _T_336 : _T_335; // @[convert.scala 46:42]
  assign _T_339 = decQ_scale[5:2]; // @[convert.scala 48:34]
  assign _T_340 = _T_339[3:3]; // @[convert.scala 49:36]
  assign _T_342 = ~ _T_339; // @[convert.scala 50:36]
  assign _T_343 = $signed(_T_342); // @[convert.scala 50:36]
  assign _T_344 = _T_340 ? $signed(_T_343) : $signed(_T_339); // @[convert.scala 50:28]
  assign _T_345 = _T_340 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_346 = ~ _T_345; // @[convert.scala 52:43]
  assign _T_350 = {_T_346,_T_345,_T_338,realFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_351 = $unsigned(_T_344); // @[Shift.scala 39:17]
  assign _T_352 = _T_351 < 4'ha; // @[Shift.scala 39:24]
  assign _T_354 = _T_350[9:8]; // @[Shift.scala 90:30]
  assign _T_355 = _T_350[7:0]; // @[Shift.scala 90:48]
  assign _T_356 = _T_355 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{1'd0}, _T_356}; // @[Shift.scala 90:39]
  assign _T_357 = _T_354 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_358 = _T_351[3]; // @[Shift.scala 12:21]
  assign _T_359 = _T_350[9]; // @[Shift.scala 12:21]
  assign _T_361 = _T_359 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_362 = {_T_361,_T_357}; // @[Cat.scala 29:58]
  assign _T_363 = _T_358 ? _T_362 : _T_350; // @[Shift.scala 91:22]
  assign _T_364 = _T_351[2:0]; // @[Shift.scala 92:77]
  assign _T_365 = _T_363[9:4]; // @[Shift.scala 90:30]
  assign _T_366 = _T_363[3:0]; // @[Shift.scala 90:48]
  assign _T_367 = _T_366 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{5'd0}, _T_367}; // @[Shift.scala 90:39]
  assign _T_368 = _T_365 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_369 = _T_364[2]; // @[Shift.scala 12:21]
  assign _T_370 = _T_363[9]; // @[Shift.scala 12:21]
  assign _T_372 = _T_370 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_373 = {_T_372,_T_368}; // @[Cat.scala 29:58]
  assign _T_374 = _T_369 ? _T_373 : _T_363; // @[Shift.scala 91:22]
  assign _T_375 = _T_364[1:0]; // @[Shift.scala 92:77]
  assign _T_376 = _T_374[9:2]; // @[Shift.scala 90:30]
  assign _T_377 = _T_374[1:0]; // @[Shift.scala 90:48]
  assign _T_378 = _T_377 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{7'd0}, _T_378}; // @[Shift.scala 90:39]
  assign _T_379 = _T_376 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_380 = _T_375[1]; // @[Shift.scala 12:21]
  assign _T_381 = _T_374[9]; // @[Shift.scala 12:21]
  assign _T_383 = _T_381 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_384 = {_T_383,_T_379}; // @[Cat.scala 29:58]
  assign _T_385 = _T_380 ? _T_384 : _T_374; // @[Shift.scala 91:22]
  assign _T_386 = _T_375[0:0]; // @[Shift.scala 92:77]
  assign _T_387 = _T_385[9:1]; // @[Shift.scala 90:30]
  assign _T_388 = _T_385[0:0]; // @[Shift.scala 90:48]
  assign _GEN_23 = {{8'd0}, _T_388}; // @[Shift.scala 90:39]
  assign _T_390 = _T_387 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_392 = _T_385[9]; // @[Shift.scala 12:21]
  assign _T_393 = {_T_392,_T_390}; // @[Cat.scala 29:58]
  assign _T_394 = _T_386 ? _T_393 : _T_385; // @[Shift.scala 91:22]
  assign _T_397 = _T_359 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_398 = _T_352 ? _T_394 : _T_397; // @[Shift.scala 39:10]
  assign _T_399 = _T_398[3]; // @[convert.scala 55:31]
  assign _T_400 = _T_398[2]; // @[convert.scala 56:31]
  assign _T_401 = _T_398[1]; // @[convert.scala 57:31]
  assign _T_402 = _T_398[0]; // @[convert.scala 58:31]
  assign _T_403 = _T_398[9:3]; // @[convert.scala 59:69]
  assign _T_404 = _T_403 != 7'h0; // @[convert.scala 59:81]
  assign _T_405 = ~ _T_404; // @[convert.scala 59:50]
  assign _T_407 = _T_403 == 7'h7f; // @[convert.scala 60:81]
  assign _T_408 = _T_399 | _T_401; // @[convert.scala 61:44]
  assign _T_409 = _T_408 | _T_402; // @[convert.scala 61:52]
  assign _T_410 = _T_400 & _T_409; // @[convert.scala 61:36]
  assign _T_411 = ~ _T_407; // @[convert.scala 62:63]
  assign _T_412 = _T_411 & _T_410; // @[convert.scala 62:103]
  assign _T_413 = _T_405 | _T_412; // @[convert.scala 62:60]
  assign _GEN_24 = {{6'd0}, _T_413}; // @[convert.scala 63:56]
  assign _T_416 = _T_403 + _GEN_24; // @[convert.scala 63:56]
  assign _T_417 = {decQ_sign,_T_416}; // @[Cat.scala 29:58]
  assign _T_419 = isZero_Z ? 8'h0 : _T_417; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 3'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_243; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 8'h80 : _T_419; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 3'h0;
    end else begin
      if (_T_202) begin
        cycleNum <= _T_219;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_186;
      end else begin
        isNaR_Z <= _T_188;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_192;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_220[4]}},_T_220};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_223) begin
      signB_Z <= _T_90;
    end
    if (_T_223) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_296) begin
      if (ready) begin
        if (_T_263) begin
          rem_Z <= _T_266;
        end else begin
          rem_Z <= _T_268;
        end
      end else begin
        if (_T_263) begin
          rem_Z <= _T_277;
        end else begin
          rem_Z <= _T_281;
        end
      end
    end
    if (_T_300) begin
      sigX_Z <= _T_311;
    end
  end
endmodule
