module PositAdder28_3(
  input         clock,
  input         reset,
  input  [27:0] io_A,
  input  [27:0] io_B,
  output [27:0] io_S
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [25:0] _T_4; // @[convert.scala 19:24]
  wire [25:0] _T_5; // @[convert.scala 19:43]
  wire [25:0] _T_6; // @[convert.scala 19:39]
  wire [15:0] _T_7; // @[LZD.scala 43:32]
  wire [7:0] _T_8; // @[LZD.scala 43:32]
  wire [3:0] _T_9; // @[LZD.scala 43:32]
  wire [1:0] _T_10; // @[LZD.scala 43:32]
  wire  _T_11; // @[LZD.scala 39:14]
  wire  _T_12; // @[LZD.scala 39:21]
  wire  _T_13; // @[LZD.scala 39:30]
  wire  _T_14; // @[LZD.scala 39:27]
  wire  _T_15; // @[LZD.scala 39:25]
  wire [1:0] _T_16; // @[Cat.scala 29:58]
  wire [1:0] _T_17; // @[LZD.scala 44:32]
  wire  _T_18; // @[LZD.scala 39:14]
  wire  _T_19; // @[LZD.scala 39:21]
  wire  _T_20; // @[LZD.scala 39:30]
  wire  _T_21; // @[LZD.scala 39:27]
  wire  _T_22; // @[LZD.scala 39:25]
  wire [1:0] _T_23; // @[Cat.scala 29:58]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[Shift.scala 12:21]
  wire  _T_26; // @[LZD.scala 49:16]
  wire  _T_27; // @[LZD.scala 49:27]
  wire  _T_28; // @[LZD.scala 49:25]
  wire  _T_29; // @[LZD.scala 49:47]
  wire  _T_30; // @[LZD.scala 49:59]
  wire  _T_31; // @[LZD.scala 49:35]
  wire [2:0] _T_33; // @[Cat.scala 29:58]
  wire [3:0] _T_34; // @[LZD.scala 44:32]
  wire [1:0] _T_35; // @[LZD.scala 43:32]
  wire  _T_36; // @[LZD.scala 39:14]
  wire  _T_37; // @[LZD.scala 39:21]
  wire  _T_38; // @[LZD.scala 39:30]
  wire  _T_39; // @[LZD.scala 39:27]
  wire  _T_40; // @[LZD.scala 39:25]
  wire [1:0] _T_41; // @[Cat.scala 29:58]
  wire [1:0] _T_42; // @[LZD.scala 44:32]
  wire  _T_43; // @[LZD.scala 39:14]
  wire  _T_44; // @[LZD.scala 39:21]
  wire  _T_45; // @[LZD.scala 39:30]
  wire  _T_46; // @[LZD.scala 39:27]
  wire  _T_47; // @[LZD.scala 39:25]
  wire [1:0] _T_48; // @[Cat.scala 29:58]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[Shift.scala 12:21]
  wire  _T_51; // @[LZD.scala 49:16]
  wire  _T_52; // @[LZD.scala 49:27]
  wire  _T_53; // @[LZD.scala 49:25]
  wire  _T_54; // @[LZD.scala 49:47]
  wire  _T_55; // @[LZD.scala 49:59]
  wire  _T_56; // @[LZD.scala 49:35]
  wire [2:0] _T_58; // @[Cat.scala 29:58]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[LZD.scala 49:16]
  wire  _T_62; // @[LZD.scala 49:27]
  wire  _T_63; // @[LZD.scala 49:25]
  wire [1:0] _T_64; // @[LZD.scala 49:47]
  wire [1:0] _T_65; // @[LZD.scala 49:59]
  wire [1:0] _T_66; // @[LZD.scala 49:35]
  wire [3:0] _T_68; // @[Cat.scala 29:58]
  wire [7:0] _T_69; // @[LZD.scala 44:32]
  wire [3:0] _T_70; // @[LZD.scala 43:32]
  wire [1:0] _T_71; // @[LZD.scala 43:32]
  wire  _T_72; // @[LZD.scala 39:14]
  wire  _T_73; // @[LZD.scala 39:21]
  wire  _T_74; // @[LZD.scala 39:30]
  wire  _T_75; // @[LZD.scala 39:27]
  wire  _T_76; // @[LZD.scala 39:25]
  wire [1:0] _T_77; // @[Cat.scala 29:58]
  wire [1:0] _T_78; // @[LZD.scala 44:32]
  wire  _T_79; // @[LZD.scala 39:14]
  wire  _T_80; // @[LZD.scala 39:21]
  wire  _T_81; // @[LZD.scala 39:30]
  wire  _T_82; // @[LZD.scala 39:27]
  wire  _T_83; // @[LZD.scala 39:25]
  wire [1:0] _T_84; // @[Cat.scala 29:58]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[Shift.scala 12:21]
  wire  _T_87; // @[LZD.scala 49:16]
  wire  _T_88; // @[LZD.scala 49:27]
  wire  _T_89; // @[LZD.scala 49:25]
  wire  _T_90; // @[LZD.scala 49:47]
  wire  _T_91; // @[LZD.scala 49:59]
  wire  _T_92; // @[LZD.scala 49:35]
  wire [2:0] _T_94; // @[Cat.scala 29:58]
  wire [3:0] _T_95; // @[LZD.scala 44:32]
  wire [1:0] _T_96; // @[LZD.scala 43:32]
  wire  _T_97; // @[LZD.scala 39:14]
  wire  _T_98; // @[LZD.scala 39:21]
  wire  _T_99; // @[LZD.scala 39:30]
  wire  _T_100; // @[LZD.scala 39:27]
  wire  _T_101; // @[LZD.scala 39:25]
  wire [1:0] _T_102; // @[Cat.scala 29:58]
  wire [1:0] _T_103; // @[LZD.scala 44:32]
  wire  _T_104; // @[LZD.scala 39:14]
  wire  _T_105; // @[LZD.scala 39:21]
  wire  _T_106; // @[LZD.scala 39:30]
  wire  _T_107; // @[LZD.scala 39:27]
  wire  _T_108; // @[LZD.scala 39:25]
  wire [1:0] _T_109; // @[Cat.scala 29:58]
  wire  _T_110; // @[Shift.scala 12:21]
  wire  _T_111; // @[Shift.scala 12:21]
  wire  _T_112; // @[LZD.scala 49:16]
  wire  _T_113; // @[LZD.scala 49:27]
  wire  _T_114; // @[LZD.scala 49:25]
  wire  _T_115; // @[LZD.scala 49:47]
  wire  _T_116; // @[LZD.scala 49:59]
  wire  _T_117; // @[LZD.scala 49:35]
  wire [2:0] _T_119; // @[Cat.scala 29:58]
  wire  _T_120; // @[Shift.scala 12:21]
  wire  _T_121; // @[Shift.scala 12:21]
  wire  _T_122; // @[LZD.scala 49:16]
  wire  _T_123; // @[LZD.scala 49:27]
  wire  _T_124; // @[LZD.scala 49:25]
  wire [1:0] _T_125; // @[LZD.scala 49:47]
  wire [1:0] _T_126; // @[LZD.scala 49:59]
  wire [1:0] _T_127; // @[LZD.scala 49:35]
  wire [3:0] _T_129; // @[Cat.scala 29:58]
  wire  _T_130; // @[Shift.scala 12:21]
  wire  _T_131; // @[Shift.scala 12:21]
  wire  _T_132; // @[LZD.scala 49:16]
  wire  _T_133; // @[LZD.scala 49:27]
  wire  _T_134; // @[LZD.scala 49:25]
  wire [2:0] _T_135; // @[LZD.scala 49:47]
  wire [2:0] _T_136; // @[LZD.scala 49:59]
  wire [2:0] _T_137; // @[LZD.scala 49:35]
  wire [4:0] _T_139; // @[Cat.scala 29:58]
  wire [9:0] _T_140; // @[LZD.scala 44:32]
  wire [7:0] _T_141; // @[LZD.scala 43:32]
  wire [3:0] _T_142; // @[LZD.scala 43:32]
  wire [1:0] _T_143; // @[LZD.scala 43:32]
  wire  _T_144; // @[LZD.scala 39:14]
  wire  _T_145; // @[LZD.scala 39:21]
  wire  _T_146; // @[LZD.scala 39:30]
  wire  _T_147; // @[LZD.scala 39:27]
  wire  _T_148; // @[LZD.scala 39:25]
  wire [1:0] _T_149; // @[Cat.scala 29:58]
  wire [1:0] _T_150; // @[LZD.scala 44:32]
  wire  _T_151; // @[LZD.scala 39:14]
  wire  _T_152; // @[LZD.scala 39:21]
  wire  _T_153; // @[LZD.scala 39:30]
  wire  _T_154; // @[LZD.scala 39:27]
  wire  _T_155; // @[LZD.scala 39:25]
  wire [1:0] _T_156; // @[Cat.scala 29:58]
  wire  _T_157; // @[Shift.scala 12:21]
  wire  _T_158; // @[Shift.scala 12:21]
  wire  _T_159; // @[LZD.scala 49:16]
  wire  _T_160; // @[LZD.scala 49:27]
  wire  _T_161; // @[LZD.scala 49:25]
  wire  _T_162; // @[LZD.scala 49:47]
  wire  _T_163; // @[LZD.scala 49:59]
  wire  _T_164; // @[LZD.scala 49:35]
  wire [2:0] _T_166; // @[Cat.scala 29:58]
  wire [3:0] _T_167; // @[LZD.scala 44:32]
  wire [1:0] _T_168; // @[LZD.scala 43:32]
  wire  _T_169; // @[LZD.scala 39:14]
  wire  _T_170; // @[LZD.scala 39:21]
  wire  _T_171; // @[LZD.scala 39:30]
  wire  _T_172; // @[LZD.scala 39:27]
  wire  _T_173; // @[LZD.scala 39:25]
  wire [1:0] _T_174; // @[Cat.scala 29:58]
  wire [1:0] _T_175; // @[LZD.scala 44:32]
  wire  _T_176; // @[LZD.scala 39:14]
  wire  _T_177; // @[LZD.scala 39:21]
  wire  _T_178; // @[LZD.scala 39:30]
  wire  _T_179; // @[LZD.scala 39:27]
  wire  _T_180; // @[LZD.scala 39:25]
  wire [1:0] _T_181; // @[Cat.scala 29:58]
  wire  _T_182; // @[Shift.scala 12:21]
  wire  _T_183; // @[Shift.scala 12:21]
  wire  _T_184; // @[LZD.scala 49:16]
  wire  _T_185; // @[LZD.scala 49:27]
  wire  _T_186; // @[LZD.scala 49:25]
  wire  _T_187; // @[LZD.scala 49:47]
  wire  _T_188; // @[LZD.scala 49:59]
  wire  _T_189; // @[LZD.scala 49:35]
  wire [2:0] _T_191; // @[Cat.scala 29:58]
  wire  _T_192; // @[Shift.scala 12:21]
  wire  _T_193; // @[Shift.scala 12:21]
  wire  _T_194; // @[LZD.scala 49:16]
  wire  _T_195; // @[LZD.scala 49:27]
  wire  _T_196; // @[LZD.scala 49:25]
  wire [1:0] _T_197; // @[LZD.scala 49:47]
  wire [1:0] _T_198; // @[LZD.scala 49:59]
  wire [1:0] _T_199; // @[LZD.scala 49:35]
  wire [3:0] _T_201; // @[Cat.scala 29:58]
  wire [1:0] _T_202; // @[LZD.scala 44:32]
  wire  _T_203; // @[LZD.scala 39:14]
  wire  _T_204; // @[LZD.scala 39:21]
  wire  _T_205; // @[LZD.scala 39:30]
  wire  _T_206; // @[LZD.scala 39:27]
  wire  _T_207; // @[LZD.scala 39:25]
  wire  _T_209; // @[Shift.scala 12:21]
  wire [2:0] _T_211; // @[Cat.scala 29:58]
  wire [2:0] _T_212; // @[LZD.scala 55:32]
  wire [2:0] _T_213; // @[LZD.scala 55:20]
  wire [3:0] _T_214; // @[Cat.scala 29:58]
  wire  _T_215; // @[Shift.scala 12:21]
  wire [3:0] _T_217; // @[LZD.scala 55:32]
  wire [3:0] _T_218; // @[LZD.scala 55:20]
  wire [4:0] _T_219; // @[Cat.scala 29:58]
  wire [4:0] _T_220; // @[convert.scala 21:22]
  wire [24:0] _T_221; // @[convert.scala 22:36]
  wire  _T_222; // @[Shift.scala 16:24]
  wire  _T_224; // @[Shift.scala 12:21]
  wire [8:0] _T_225; // @[Shift.scala 64:52]
  wire [24:0] _T_227; // @[Cat.scala 29:58]
  wire [24:0] _T_228; // @[Shift.scala 64:27]
  wire [3:0] _T_229; // @[Shift.scala 66:70]
  wire  _T_230; // @[Shift.scala 12:21]
  wire [16:0] _T_231; // @[Shift.scala 64:52]
  wire [24:0] _T_233; // @[Cat.scala 29:58]
  wire [24:0] _T_234; // @[Shift.scala 64:27]
  wire [2:0] _T_235; // @[Shift.scala 66:70]
  wire  _T_236; // @[Shift.scala 12:21]
  wire [20:0] _T_237; // @[Shift.scala 64:52]
  wire [24:0] _T_239; // @[Cat.scala 29:58]
  wire [24:0] _T_240; // @[Shift.scala 64:27]
  wire [1:0] _T_241; // @[Shift.scala 66:70]
  wire  _T_242; // @[Shift.scala 12:21]
  wire [22:0] _T_243; // @[Shift.scala 64:52]
  wire [24:0] _T_245; // @[Cat.scala 29:58]
  wire [24:0] _T_246; // @[Shift.scala 64:27]
  wire  _T_247; // @[Shift.scala 66:70]
  wire [23:0] _T_249; // @[Shift.scala 64:52]
  wire [24:0] _T_250; // @[Cat.scala 29:58]
  wire [24:0] _T_251; // @[Shift.scala 64:27]
  wire [24:0] _T_252; // @[Shift.scala 16:10]
  wire [2:0] _T_253; // @[convert.scala 23:34]
  wire [21:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_255; // @[convert.scala 25:26]
  wire [4:0] _T_257; // @[convert.scala 25:42]
  wire [2:0] _T_260; // @[convert.scala 26:67]
  wire [2:0] _T_261; // @[convert.scala 26:51]
  wire [8:0] _T_262; // @[Cat.scala 29:58]
  wire [26:0] _T_264; // @[convert.scala 29:56]
  wire  _T_265; // @[convert.scala 29:60]
  wire  _T_266; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_269; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [8:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_278; // @[convert.scala 18:24]
  wire  _T_279; // @[convert.scala 18:40]
  wire  _T_280; // @[convert.scala 18:36]
  wire [25:0] _T_281; // @[convert.scala 19:24]
  wire [25:0] _T_282; // @[convert.scala 19:43]
  wire [25:0] _T_283; // @[convert.scala 19:39]
  wire [15:0] _T_284; // @[LZD.scala 43:32]
  wire [7:0] _T_285; // @[LZD.scala 43:32]
  wire [3:0] _T_286; // @[LZD.scala 43:32]
  wire [1:0] _T_287; // @[LZD.scala 43:32]
  wire  _T_288; // @[LZD.scala 39:14]
  wire  _T_289; // @[LZD.scala 39:21]
  wire  _T_290; // @[LZD.scala 39:30]
  wire  _T_291; // @[LZD.scala 39:27]
  wire  _T_292; // @[LZD.scala 39:25]
  wire [1:0] _T_293; // @[Cat.scala 29:58]
  wire [1:0] _T_294; // @[LZD.scala 44:32]
  wire  _T_295; // @[LZD.scala 39:14]
  wire  _T_296; // @[LZD.scala 39:21]
  wire  _T_297; // @[LZD.scala 39:30]
  wire  _T_298; // @[LZD.scala 39:27]
  wire  _T_299; // @[LZD.scala 39:25]
  wire [1:0] _T_300; // @[Cat.scala 29:58]
  wire  _T_301; // @[Shift.scala 12:21]
  wire  _T_302; // @[Shift.scala 12:21]
  wire  _T_303; // @[LZD.scala 49:16]
  wire  _T_304; // @[LZD.scala 49:27]
  wire  _T_305; // @[LZD.scala 49:25]
  wire  _T_306; // @[LZD.scala 49:47]
  wire  _T_307; // @[LZD.scala 49:59]
  wire  _T_308; // @[LZD.scala 49:35]
  wire [2:0] _T_310; // @[Cat.scala 29:58]
  wire [3:0] _T_311; // @[LZD.scala 44:32]
  wire [1:0] _T_312; // @[LZD.scala 43:32]
  wire  _T_313; // @[LZD.scala 39:14]
  wire  _T_314; // @[LZD.scala 39:21]
  wire  _T_315; // @[LZD.scala 39:30]
  wire  _T_316; // @[LZD.scala 39:27]
  wire  _T_317; // @[LZD.scala 39:25]
  wire [1:0] _T_318; // @[Cat.scala 29:58]
  wire [1:0] _T_319; // @[LZD.scala 44:32]
  wire  _T_320; // @[LZD.scala 39:14]
  wire  _T_321; // @[LZD.scala 39:21]
  wire  _T_322; // @[LZD.scala 39:30]
  wire  _T_323; // @[LZD.scala 39:27]
  wire  _T_324; // @[LZD.scala 39:25]
  wire [1:0] _T_325; // @[Cat.scala 29:58]
  wire  _T_326; // @[Shift.scala 12:21]
  wire  _T_327; // @[Shift.scala 12:21]
  wire  _T_328; // @[LZD.scala 49:16]
  wire  _T_329; // @[LZD.scala 49:27]
  wire  _T_330; // @[LZD.scala 49:25]
  wire  _T_331; // @[LZD.scala 49:47]
  wire  _T_332; // @[LZD.scala 49:59]
  wire  _T_333; // @[LZD.scala 49:35]
  wire [2:0] _T_335; // @[Cat.scala 29:58]
  wire  _T_336; // @[Shift.scala 12:21]
  wire  _T_337; // @[Shift.scala 12:21]
  wire  _T_338; // @[LZD.scala 49:16]
  wire  _T_339; // @[LZD.scala 49:27]
  wire  _T_340; // @[LZD.scala 49:25]
  wire [1:0] _T_341; // @[LZD.scala 49:47]
  wire [1:0] _T_342; // @[LZD.scala 49:59]
  wire [1:0] _T_343; // @[LZD.scala 49:35]
  wire [3:0] _T_345; // @[Cat.scala 29:58]
  wire [7:0] _T_346; // @[LZD.scala 44:32]
  wire [3:0] _T_347; // @[LZD.scala 43:32]
  wire [1:0] _T_348; // @[LZD.scala 43:32]
  wire  _T_349; // @[LZD.scala 39:14]
  wire  _T_350; // @[LZD.scala 39:21]
  wire  _T_351; // @[LZD.scala 39:30]
  wire  _T_352; // @[LZD.scala 39:27]
  wire  _T_353; // @[LZD.scala 39:25]
  wire [1:0] _T_354; // @[Cat.scala 29:58]
  wire [1:0] _T_355; // @[LZD.scala 44:32]
  wire  _T_356; // @[LZD.scala 39:14]
  wire  _T_357; // @[LZD.scala 39:21]
  wire  _T_358; // @[LZD.scala 39:30]
  wire  _T_359; // @[LZD.scala 39:27]
  wire  _T_360; // @[LZD.scala 39:25]
  wire [1:0] _T_361; // @[Cat.scala 29:58]
  wire  _T_362; // @[Shift.scala 12:21]
  wire  _T_363; // @[Shift.scala 12:21]
  wire  _T_364; // @[LZD.scala 49:16]
  wire  _T_365; // @[LZD.scala 49:27]
  wire  _T_366; // @[LZD.scala 49:25]
  wire  _T_367; // @[LZD.scala 49:47]
  wire  _T_368; // @[LZD.scala 49:59]
  wire  _T_369; // @[LZD.scala 49:35]
  wire [2:0] _T_371; // @[Cat.scala 29:58]
  wire [3:0] _T_372; // @[LZD.scala 44:32]
  wire [1:0] _T_373; // @[LZD.scala 43:32]
  wire  _T_374; // @[LZD.scala 39:14]
  wire  _T_375; // @[LZD.scala 39:21]
  wire  _T_376; // @[LZD.scala 39:30]
  wire  _T_377; // @[LZD.scala 39:27]
  wire  _T_378; // @[LZD.scala 39:25]
  wire [1:0] _T_379; // @[Cat.scala 29:58]
  wire [1:0] _T_380; // @[LZD.scala 44:32]
  wire  _T_381; // @[LZD.scala 39:14]
  wire  _T_382; // @[LZD.scala 39:21]
  wire  _T_383; // @[LZD.scala 39:30]
  wire  _T_384; // @[LZD.scala 39:27]
  wire  _T_385; // @[LZD.scala 39:25]
  wire [1:0] _T_386; // @[Cat.scala 29:58]
  wire  _T_387; // @[Shift.scala 12:21]
  wire  _T_388; // @[Shift.scala 12:21]
  wire  _T_389; // @[LZD.scala 49:16]
  wire  _T_390; // @[LZD.scala 49:27]
  wire  _T_391; // @[LZD.scala 49:25]
  wire  _T_392; // @[LZD.scala 49:47]
  wire  _T_393; // @[LZD.scala 49:59]
  wire  _T_394; // @[LZD.scala 49:35]
  wire [2:0] _T_396; // @[Cat.scala 29:58]
  wire  _T_397; // @[Shift.scala 12:21]
  wire  _T_398; // @[Shift.scala 12:21]
  wire  _T_399; // @[LZD.scala 49:16]
  wire  _T_400; // @[LZD.scala 49:27]
  wire  _T_401; // @[LZD.scala 49:25]
  wire [1:0] _T_402; // @[LZD.scala 49:47]
  wire [1:0] _T_403; // @[LZD.scala 49:59]
  wire [1:0] _T_404; // @[LZD.scala 49:35]
  wire [3:0] _T_406; // @[Cat.scala 29:58]
  wire  _T_407; // @[Shift.scala 12:21]
  wire  _T_408; // @[Shift.scala 12:21]
  wire  _T_409; // @[LZD.scala 49:16]
  wire  _T_410; // @[LZD.scala 49:27]
  wire  _T_411; // @[LZD.scala 49:25]
  wire [2:0] _T_412; // @[LZD.scala 49:47]
  wire [2:0] _T_413; // @[LZD.scala 49:59]
  wire [2:0] _T_414; // @[LZD.scala 49:35]
  wire [4:0] _T_416; // @[Cat.scala 29:58]
  wire [9:0] _T_417; // @[LZD.scala 44:32]
  wire [7:0] _T_418; // @[LZD.scala 43:32]
  wire [3:0] _T_419; // @[LZD.scala 43:32]
  wire [1:0] _T_420; // @[LZD.scala 43:32]
  wire  _T_421; // @[LZD.scala 39:14]
  wire  _T_422; // @[LZD.scala 39:21]
  wire  _T_423; // @[LZD.scala 39:30]
  wire  _T_424; // @[LZD.scala 39:27]
  wire  _T_425; // @[LZD.scala 39:25]
  wire [1:0] _T_426; // @[Cat.scala 29:58]
  wire [1:0] _T_427; // @[LZD.scala 44:32]
  wire  _T_428; // @[LZD.scala 39:14]
  wire  _T_429; // @[LZD.scala 39:21]
  wire  _T_430; // @[LZD.scala 39:30]
  wire  _T_431; // @[LZD.scala 39:27]
  wire  _T_432; // @[LZD.scala 39:25]
  wire [1:0] _T_433; // @[Cat.scala 29:58]
  wire  _T_434; // @[Shift.scala 12:21]
  wire  _T_435; // @[Shift.scala 12:21]
  wire  _T_436; // @[LZD.scala 49:16]
  wire  _T_437; // @[LZD.scala 49:27]
  wire  _T_438; // @[LZD.scala 49:25]
  wire  _T_439; // @[LZD.scala 49:47]
  wire  _T_440; // @[LZD.scala 49:59]
  wire  _T_441; // @[LZD.scala 49:35]
  wire [2:0] _T_443; // @[Cat.scala 29:58]
  wire [3:0] _T_444; // @[LZD.scala 44:32]
  wire [1:0] _T_445; // @[LZD.scala 43:32]
  wire  _T_446; // @[LZD.scala 39:14]
  wire  _T_447; // @[LZD.scala 39:21]
  wire  _T_448; // @[LZD.scala 39:30]
  wire  _T_449; // @[LZD.scala 39:27]
  wire  _T_450; // @[LZD.scala 39:25]
  wire [1:0] _T_451; // @[Cat.scala 29:58]
  wire [1:0] _T_452; // @[LZD.scala 44:32]
  wire  _T_453; // @[LZD.scala 39:14]
  wire  _T_454; // @[LZD.scala 39:21]
  wire  _T_455; // @[LZD.scala 39:30]
  wire  _T_456; // @[LZD.scala 39:27]
  wire  _T_457; // @[LZD.scala 39:25]
  wire [1:0] _T_458; // @[Cat.scala 29:58]
  wire  _T_459; // @[Shift.scala 12:21]
  wire  _T_460; // @[Shift.scala 12:21]
  wire  _T_461; // @[LZD.scala 49:16]
  wire  _T_462; // @[LZD.scala 49:27]
  wire  _T_463; // @[LZD.scala 49:25]
  wire  _T_464; // @[LZD.scala 49:47]
  wire  _T_465; // @[LZD.scala 49:59]
  wire  _T_466; // @[LZD.scala 49:35]
  wire [2:0] _T_468; // @[Cat.scala 29:58]
  wire  _T_469; // @[Shift.scala 12:21]
  wire  _T_470; // @[Shift.scala 12:21]
  wire  _T_471; // @[LZD.scala 49:16]
  wire  _T_472; // @[LZD.scala 49:27]
  wire  _T_473; // @[LZD.scala 49:25]
  wire [1:0] _T_474; // @[LZD.scala 49:47]
  wire [1:0] _T_475; // @[LZD.scala 49:59]
  wire [1:0] _T_476; // @[LZD.scala 49:35]
  wire [3:0] _T_478; // @[Cat.scala 29:58]
  wire [1:0] _T_479; // @[LZD.scala 44:32]
  wire  _T_480; // @[LZD.scala 39:14]
  wire  _T_481; // @[LZD.scala 39:21]
  wire  _T_482; // @[LZD.scala 39:30]
  wire  _T_483; // @[LZD.scala 39:27]
  wire  _T_484; // @[LZD.scala 39:25]
  wire  _T_486; // @[Shift.scala 12:21]
  wire [2:0] _T_488; // @[Cat.scala 29:58]
  wire [2:0] _T_489; // @[LZD.scala 55:32]
  wire [2:0] _T_490; // @[LZD.scala 55:20]
  wire [3:0] _T_491; // @[Cat.scala 29:58]
  wire  _T_492; // @[Shift.scala 12:21]
  wire [3:0] _T_494; // @[LZD.scala 55:32]
  wire [3:0] _T_495; // @[LZD.scala 55:20]
  wire [4:0] _T_496; // @[Cat.scala 29:58]
  wire [4:0] _T_497; // @[convert.scala 21:22]
  wire [24:0] _T_498; // @[convert.scala 22:36]
  wire  _T_499; // @[Shift.scala 16:24]
  wire  _T_501; // @[Shift.scala 12:21]
  wire [8:0] _T_502; // @[Shift.scala 64:52]
  wire [24:0] _T_504; // @[Cat.scala 29:58]
  wire [24:0] _T_505; // @[Shift.scala 64:27]
  wire [3:0] _T_506; // @[Shift.scala 66:70]
  wire  _T_507; // @[Shift.scala 12:21]
  wire [16:0] _T_508; // @[Shift.scala 64:52]
  wire [24:0] _T_510; // @[Cat.scala 29:58]
  wire [24:0] _T_511; // @[Shift.scala 64:27]
  wire [2:0] _T_512; // @[Shift.scala 66:70]
  wire  _T_513; // @[Shift.scala 12:21]
  wire [20:0] _T_514; // @[Shift.scala 64:52]
  wire [24:0] _T_516; // @[Cat.scala 29:58]
  wire [24:0] _T_517; // @[Shift.scala 64:27]
  wire [1:0] _T_518; // @[Shift.scala 66:70]
  wire  _T_519; // @[Shift.scala 12:21]
  wire [22:0] _T_520; // @[Shift.scala 64:52]
  wire [24:0] _T_522; // @[Cat.scala 29:58]
  wire [24:0] _T_523; // @[Shift.scala 64:27]
  wire  _T_524; // @[Shift.scala 66:70]
  wire [23:0] _T_526; // @[Shift.scala 64:52]
  wire [24:0] _T_527; // @[Cat.scala 29:58]
  wire [24:0] _T_528; // @[Shift.scala 64:27]
  wire [24:0] _T_529; // @[Shift.scala 16:10]
  wire [2:0] _T_530; // @[convert.scala 23:34]
  wire [21:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_532; // @[convert.scala 25:26]
  wire [4:0] _T_534; // @[convert.scala 25:42]
  wire [2:0] _T_537; // @[convert.scala 26:67]
  wire [2:0] _T_538; // @[convert.scala 26:51]
  wire [8:0] _T_539; // @[Cat.scala 29:58]
  wire [26:0] _T_541; // @[convert.scala 29:56]
  wire  _T_542; // @[convert.scala 29:60]
  wire  _T_543; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_546; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [8:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[PositAdder.scala 24:32]
  wire  greaterSign; // @[PositAdder.scala 25:24]
  wire  smallerSign; // @[PositAdder.scala 26:24]
  wire [8:0] greaterExp; // @[PositAdder.scala 27:24]
  wire [8:0] smallerExp; // @[PositAdder.scala 28:24]
  wire [21:0] greaterFrac; // @[PositAdder.scala 29:24]
  wire [21:0] smallerFrac; // @[PositAdder.scala 30:24]
  wire [8:0] _T_555; // @[PositAdder.scala 31:32]
  wire [8:0] scale_diff; // @[PositAdder.scala 31:32]
  wire  _T_556; // @[PositAdder.scala 32:38]
  wire [23:0] greaterSig; // @[Cat.scala 29:58]
  wire  _T_558; // @[PositAdder.scala 33:38]
  wire [26:0] _T_561; // @[Cat.scala 29:58]
  wire [8:0] _T_562; // @[PositAdder.scala 34:68]
  wire  _T_563; // @[Shift.scala 39:24]
  wire [4:0] _T_564; // @[Shift.scala 40:44]
  wire [10:0] _T_565; // @[Shift.scala 90:30]
  wire [15:0] _T_566; // @[Shift.scala 90:48]
  wire  _T_567; // @[Shift.scala 90:57]
  wire [10:0] _GEN_0; // @[Shift.scala 90:39]
  wire [10:0] _T_568; // @[Shift.scala 90:39]
  wire  _T_569; // @[Shift.scala 12:21]
  wire  _T_570; // @[Shift.scala 12:21]
  wire [15:0] _T_572; // @[Bitwise.scala 71:12]
  wire [26:0] _T_573; // @[Cat.scala 29:58]
  wire [26:0] _T_574; // @[Shift.scala 91:22]
  wire [3:0] _T_575; // @[Shift.scala 92:77]
  wire [18:0] _T_576; // @[Shift.scala 90:30]
  wire [7:0] _T_577; // @[Shift.scala 90:48]
  wire  _T_578; // @[Shift.scala 90:57]
  wire [18:0] _GEN_1; // @[Shift.scala 90:39]
  wire [18:0] _T_579; // @[Shift.scala 90:39]
  wire  _T_580; // @[Shift.scala 12:21]
  wire  _T_581; // @[Shift.scala 12:21]
  wire [7:0] _T_583; // @[Bitwise.scala 71:12]
  wire [26:0] _T_584; // @[Cat.scala 29:58]
  wire [26:0] _T_585; // @[Shift.scala 91:22]
  wire [2:0] _T_586; // @[Shift.scala 92:77]
  wire [22:0] _T_587; // @[Shift.scala 90:30]
  wire [3:0] _T_588; // @[Shift.scala 90:48]
  wire  _T_589; // @[Shift.scala 90:57]
  wire [22:0] _GEN_2; // @[Shift.scala 90:39]
  wire [22:0] _T_590; // @[Shift.scala 90:39]
  wire  _T_591; // @[Shift.scala 12:21]
  wire  _T_592; // @[Shift.scala 12:21]
  wire [3:0] _T_594; // @[Bitwise.scala 71:12]
  wire [26:0] _T_595; // @[Cat.scala 29:58]
  wire [26:0] _T_596; // @[Shift.scala 91:22]
  wire [1:0] _T_597; // @[Shift.scala 92:77]
  wire [24:0] _T_598; // @[Shift.scala 90:30]
  wire [1:0] _T_599; // @[Shift.scala 90:48]
  wire  _T_600; // @[Shift.scala 90:57]
  wire [24:0] _GEN_3; // @[Shift.scala 90:39]
  wire [24:0] _T_601; // @[Shift.scala 90:39]
  wire  _T_602; // @[Shift.scala 12:21]
  wire  _T_603; // @[Shift.scala 12:21]
  wire [1:0] _T_605; // @[Bitwise.scala 71:12]
  wire [26:0] _T_606; // @[Cat.scala 29:58]
  wire [26:0] _T_607; // @[Shift.scala 91:22]
  wire  _T_608; // @[Shift.scala 92:77]
  wire [25:0] _T_609; // @[Shift.scala 90:30]
  wire  _T_610; // @[Shift.scala 90:48]
  wire [25:0] _GEN_4; // @[Shift.scala 90:39]
  wire [25:0] _T_612; // @[Shift.scala 90:39]
  wire  _T_614; // @[Shift.scala 12:21]
  wire [26:0] _T_615; // @[Cat.scala 29:58]
  wire [26:0] _T_616; // @[Shift.scala 91:22]
  wire [26:0] _T_619; // @[Bitwise.scala 71:12]
  wire [26:0] smallerSig; // @[Shift.scala 39:10]
  wire [23:0] _T_620; // @[PositAdder.scala 35:45]
  wire [24:0] rawSumSig; // @[PositAdder.scala 35:32]
  wire  _T_621; // @[PositAdder.scala 36:31]
  wire  _T_622; // @[PositAdder.scala 36:59]
  wire  sumSign; // @[PositAdder.scala 36:43]
  wire [23:0] _T_623; // @[PositAdder.scala 37:48]
  wire [2:0] _T_624; // @[PositAdder.scala 37:63]
  wire [27:0] signSumSig; // @[Cat.scala 29:58]
  wire [26:0] _T_626; // @[PositAdder.scala 39:31]
  wire [26:0] _T_627; // @[PositAdder.scala 39:66]
  wire [26:0] sumXor; // @[PositAdder.scala 39:49]
  wire [15:0] _T_628; // @[LZD.scala 43:32]
  wire [7:0] _T_629; // @[LZD.scala 43:32]
  wire [3:0] _T_630; // @[LZD.scala 43:32]
  wire [1:0] _T_631; // @[LZD.scala 43:32]
  wire  _T_632; // @[LZD.scala 39:14]
  wire  _T_633; // @[LZD.scala 39:21]
  wire  _T_634; // @[LZD.scala 39:30]
  wire  _T_635; // @[LZD.scala 39:27]
  wire  _T_636; // @[LZD.scala 39:25]
  wire [1:0] _T_637; // @[Cat.scala 29:58]
  wire [1:0] _T_638; // @[LZD.scala 44:32]
  wire  _T_639; // @[LZD.scala 39:14]
  wire  _T_640; // @[LZD.scala 39:21]
  wire  _T_641; // @[LZD.scala 39:30]
  wire  _T_642; // @[LZD.scala 39:27]
  wire  _T_643; // @[LZD.scala 39:25]
  wire [1:0] _T_644; // @[Cat.scala 29:58]
  wire  _T_645; // @[Shift.scala 12:21]
  wire  _T_646; // @[Shift.scala 12:21]
  wire  _T_647; // @[LZD.scala 49:16]
  wire  _T_648; // @[LZD.scala 49:27]
  wire  _T_649; // @[LZD.scala 49:25]
  wire  _T_650; // @[LZD.scala 49:47]
  wire  _T_651; // @[LZD.scala 49:59]
  wire  _T_652; // @[LZD.scala 49:35]
  wire [2:0] _T_654; // @[Cat.scala 29:58]
  wire [3:0] _T_655; // @[LZD.scala 44:32]
  wire [1:0] _T_656; // @[LZD.scala 43:32]
  wire  _T_657; // @[LZD.scala 39:14]
  wire  _T_658; // @[LZD.scala 39:21]
  wire  _T_659; // @[LZD.scala 39:30]
  wire  _T_660; // @[LZD.scala 39:27]
  wire  _T_661; // @[LZD.scala 39:25]
  wire [1:0] _T_662; // @[Cat.scala 29:58]
  wire [1:0] _T_663; // @[LZD.scala 44:32]
  wire  _T_664; // @[LZD.scala 39:14]
  wire  _T_665; // @[LZD.scala 39:21]
  wire  _T_666; // @[LZD.scala 39:30]
  wire  _T_667; // @[LZD.scala 39:27]
  wire  _T_668; // @[LZD.scala 39:25]
  wire [1:0] _T_669; // @[Cat.scala 29:58]
  wire  _T_670; // @[Shift.scala 12:21]
  wire  _T_671; // @[Shift.scala 12:21]
  wire  _T_672; // @[LZD.scala 49:16]
  wire  _T_673; // @[LZD.scala 49:27]
  wire  _T_674; // @[LZD.scala 49:25]
  wire  _T_675; // @[LZD.scala 49:47]
  wire  _T_676; // @[LZD.scala 49:59]
  wire  _T_677; // @[LZD.scala 49:35]
  wire [2:0] _T_679; // @[Cat.scala 29:58]
  wire  _T_680; // @[Shift.scala 12:21]
  wire  _T_681; // @[Shift.scala 12:21]
  wire  _T_682; // @[LZD.scala 49:16]
  wire  _T_683; // @[LZD.scala 49:27]
  wire  _T_684; // @[LZD.scala 49:25]
  wire [1:0] _T_685; // @[LZD.scala 49:47]
  wire [1:0] _T_686; // @[LZD.scala 49:59]
  wire [1:0] _T_687; // @[LZD.scala 49:35]
  wire [3:0] _T_689; // @[Cat.scala 29:58]
  wire [7:0] _T_690; // @[LZD.scala 44:32]
  wire [3:0] _T_691; // @[LZD.scala 43:32]
  wire [1:0] _T_692; // @[LZD.scala 43:32]
  wire  _T_693; // @[LZD.scala 39:14]
  wire  _T_694; // @[LZD.scala 39:21]
  wire  _T_695; // @[LZD.scala 39:30]
  wire  _T_696; // @[LZD.scala 39:27]
  wire  _T_697; // @[LZD.scala 39:25]
  wire [1:0] _T_698; // @[Cat.scala 29:58]
  wire [1:0] _T_699; // @[LZD.scala 44:32]
  wire  _T_700; // @[LZD.scala 39:14]
  wire  _T_701; // @[LZD.scala 39:21]
  wire  _T_702; // @[LZD.scala 39:30]
  wire  _T_703; // @[LZD.scala 39:27]
  wire  _T_704; // @[LZD.scala 39:25]
  wire [1:0] _T_705; // @[Cat.scala 29:58]
  wire  _T_706; // @[Shift.scala 12:21]
  wire  _T_707; // @[Shift.scala 12:21]
  wire  _T_708; // @[LZD.scala 49:16]
  wire  _T_709; // @[LZD.scala 49:27]
  wire  _T_710; // @[LZD.scala 49:25]
  wire  _T_711; // @[LZD.scala 49:47]
  wire  _T_712; // @[LZD.scala 49:59]
  wire  _T_713; // @[LZD.scala 49:35]
  wire [2:0] _T_715; // @[Cat.scala 29:58]
  wire [3:0] _T_716; // @[LZD.scala 44:32]
  wire [1:0] _T_717; // @[LZD.scala 43:32]
  wire  _T_718; // @[LZD.scala 39:14]
  wire  _T_719; // @[LZD.scala 39:21]
  wire  _T_720; // @[LZD.scala 39:30]
  wire  _T_721; // @[LZD.scala 39:27]
  wire  _T_722; // @[LZD.scala 39:25]
  wire [1:0] _T_723; // @[Cat.scala 29:58]
  wire [1:0] _T_724; // @[LZD.scala 44:32]
  wire  _T_725; // @[LZD.scala 39:14]
  wire  _T_726; // @[LZD.scala 39:21]
  wire  _T_727; // @[LZD.scala 39:30]
  wire  _T_728; // @[LZD.scala 39:27]
  wire  _T_729; // @[LZD.scala 39:25]
  wire [1:0] _T_730; // @[Cat.scala 29:58]
  wire  _T_731; // @[Shift.scala 12:21]
  wire  _T_732; // @[Shift.scala 12:21]
  wire  _T_733; // @[LZD.scala 49:16]
  wire  _T_734; // @[LZD.scala 49:27]
  wire  _T_735; // @[LZD.scala 49:25]
  wire  _T_736; // @[LZD.scala 49:47]
  wire  _T_737; // @[LZD.scala 49:59]
  wire  _T_738; // @[LZD.scala 49:35]
  wire [2:0] _T_740; // @[Cat.scala 29:58]
  wire  _T_741; // @[Shift.scala 12:21]
  wire  _T_742; // @[Shift.scala 12:21]
  wire  _T_743; // @[LZD.scala 49:16]
  wire  _T_744; // @[LZD.scala 49:27]
  wire  _T_745; // @[LZD.scala 49:25]
  wire [1:0] _T_746; // @[LZD.scala 49:47]
  wire [1:0] _T_747; // @[LZD.scala 49:59]
  wire [1:0] _T_748; // @[LZD.scala 49:35]
  wire [3:0] _T_750; // @[Cat.scala 29:58]
  wire  _T_751; // @[Shift.scala 12:21]
  wire  _T_752; // @[Shift.scala 12:21]
  wire  _T_753; // @[LZD.scala 49:16]
  wire  _T_754; // @[LZD.scala 49:27]
  wire  _T_755; // @[LZD.scala 49:25]
  wire [2:0] _T_756; // @[LZD.scala 49:47]
  wire [2:0] _T_757; // @[LZD.scala 49:59]
  wire [2:0] _T_758; // @[LZD.scala 49:35]
  wire [4:0] _T_760; // @[Cat.scala 29:58]
  wire [10:0] _T_761; // @[LZD.scala 44:32]
  wire [7:0] _T_762; // @[LZD.scala 43:32]
  wire [3:0] _T_763; // @[LZD.scala 43:32]
  wire [1:0] _T_764; // @[LZD.scala 43:32]
  wire  _T_765; // @[LZD.scala 39:14]
  wire  _T_766; // @[LZD.scala 39:21]
  wire  _T_767; // @[LZD.scala 39:30]
  wire  _T_768; // @[LZD.scala 39:27]
  wire  _T_769; // @[LZD.scala 39:25]
  wire [1:0] _T_770; // @[Cat.scala 29:58]
  wire [1:0] _T_771; // @[LZD.scala 44:32]
  wire  _T_772; // @[LZD.scala 39:14]
  wire  _T_773; // @[LZD.scala 39:21]
  wire  _T_774; // @[LZD.scala 39:30]
  wire  _T_775; // @[LZD.scala 39:27]
  wire  _T_776; // @[LZD.scala 39:25]
  wire [1:0] _T_777; // @[Cat.scala 29:58]
  wire  _T_778; // @[Shift.scala 12:21]
  wire  _T_779; // @[Shift.scala 12:21]
  wire  _T_780; // @[LZD.scala 49:16]
  wire  _T_781; // @[LZD.scala 49:27]
  wire  _T_782; // @[LZD.scala 49:25]
  wire  _T_783; // @[LZD.scala 49:47]
  wire  _T_784; // @[LZD.scala 49:59]
  wire  _T_785; // @[LZD.scala 49:35]
  wire [2:0] _T_787; // @[Cat.scala 29:58]
  wire [3:0] _T_788; // @[LZD.scala 44:32]
  wire [1:0] _T_789; // @[LZD.scala 43:32]
  wire  _T_790; // @[LZD.scala 39:14]
  wire  _T_791; // @[LZD.scala 39:21]
  wire  _T_792; // @[LZD.scala 39:30]
  wire  _T_793; // @[LZD.scala 39:27]
  wire  _T_794; // @[LZD.scala 39:25]
  wire [1:0] _T_795; // @[Cat.scala 29:58]
  wire [1:0] _T_796; // @[LZD.scala 44:32]
  wire  _T_797; // @[LZD.scala 39:14]
  wire  _T_798; // @[LZD.scala 39:21]
  wire  _T_799; // @[LZD.scala 39:30]
  wire  _T_800; // @[LZD.scala 39:27]
  wire  _T_801; // @[LZD.scala 39:25]
  wire [1:0] _T_802; // @[Cat.scala 29:58]
  wire  _T_803; // @[Shift.scala 12:21]
  wire  _T_804; // @[Shift.scala 12:21]
  wire  _T_805; // @[LZD.scala 49:16]
  wire  _T_806; // @[LZD.scala 49:27]
  wire  _T_807; // @[LZD.scala 49:25]
  wire  _T_808; // @[LZD.scala 49:47]
  wire  _T_809; // @[LZD.scala 49:59]
  wire  _T_810; // @[LZD.scala 49:35]
  wire [2:0] _T_812; // @[Cat.scala 29:58]
  wire  _T_813; // @[Shift.scala 12:21]
  wire  _T_814; // @[Shift.scala 12:21]
  wire  _T_815; // @[LZD.scala 49:16]
  wire  _T_816; // @[LZD.scala 49:27]
  wire  _T_817; // @[LZD.scala 49:25]
  wire [1:0] _T_818; // @[LZD.scala 49:47]
  wire [1:0] _T_819; // @[LZD.scala 49:59]
  wire [1:0] _T_820; // @[LZD.scala 49:35]
  wire [3:0] _T_822; // @[Cat.scala 29:58]
  wire [2:0] _T_823; // @[LZD.scala 44:32]
  wire [1:0] _T_824; // @[LZD.scala 43:32]
  wire  _T_825; // @[LZD.scala 39:14]
  wire  _T_826; // @[LZD.scala 39:21]
  wire  _T_827; // @[LZD.scala 39:30]
  wire  _T_828; // @[LZD.scala 39:27]
  wire  _T_829; // @[LZD.scala 39:25]
  wire [1:0] _T_830; // @[Cat.scala 29:58]
  wire  _T_831; // @[LZD.scala 44:32]
  wire  _T_833; // @[Shift.scala 12:21]
  wire  _T_835; // @[LZD.scala 55:32]
  wire  _T_836; // @[LZD.scala 55:20]
  wire  _T_838; // @[Shift.scala 12:21]
  wire [2:0] _T_840; // @[Cat.scala 29:58]
  wire [2:0] _T_841; // @[LZD.scala 55:32]
  wire [2:0] _T_842; // @[LZD.scala 55:20]
  wire [3:0] _T_843; // @[Cat.scala 29:58]
  wire  _T_844; // @[Shift.scala 12:21]
  wire [3:0] _T_846; // @[LZD.scala 55:32]
  wire [3:0] _T_847; // @[LZD.scala 55:20]
  wire [4:0] sumLZD; // @[Cat.scala 29:58]
  wire [5:0] _T_848; // @[Cat.scala 29:58]
  wire [5:0] _T_849; // @[PositAdder.scala 41:38]
  wire [5:0] _T_851; // @[PositAdder.scala 41:45]
  wire [5:0] scaleBias; // @[PositAdder.scala 41:45]
  wire [8:0] _GEN_5; // @[PositAdder.scala 42:32]
  wire [9:0] sumScale; // @[PositAdder.scala 42:32]
  wire  overflow; // @[PositAdder.scala 43:30]
  wire [4:0] normalShift; // @[PositAdder.scala 44:22]
  wire [25:0] _T_852; // @[PositAdder.scala 45:36]
  wire  _T_853; // @[Shift.scala 16:24]
  wire  _T_855; // @[Shift.scala 12:21]
  wire [9:0] _T_856; // @[Shift.scala 64:52]
  wire [25:0] _T_858; // @[Cat.scala 29:58]
  wire [25:0] _T_859; // @[Shift.scala 64:27]
  wire [3:0] _T_860; // @[Shift.scala 66:70]
  wire  _T_861; // @[Shift.scala 12:21]
  wire [17:0] _T_862; // @[Shift.scala 64:52]
  wire [25:0] _T_864; // @[Cat.scala 29:58]
  wire [25:0] _T_865; // @[Shift.scala 64:27]
  wire [2:0] _T_866; // @[Shift.scala 66:70]
  wire  _T_867; // @[Shift.scala 12:21]
  wire [21:0] _T_868; // @[Shift.scala 64:52]
  wire [25:0] _T_870; // @[Cat.scala 29:58]
  wire [25:0] _T_871; // @[Shift.scala 64:27]
  wire [1:0] _T_872; // @[Shift.scala 66:70]
  wire  _T_873; // @[Shift.scala 12:21]
  wire [23:0] _T_874; // @[Shift.scala 64:52]
  wire [25:0] _T_876; // @[Cat.scala 29:58]
  wire [25:0] _T_877; // @[Shift.scala 64:27]
  wire  _T_878; // @[Shift.scala 66:70]
  wire [24:0] _T_880; // @[Shift.scala 64:52]
  wire [25:0] _T_881; // @[Cat.scala 29:58]
  wire [25:0] _T_882; // @[Shift.scala 64:27]
  wire [25:0] shiftSig; // @[Shift.scala 16:10]
  wire [9:0] _T_883; // @[PositAdder.scala 50:24]
  wire [21:0] decS_fraction; // @[PositAdder.scala 51:34]
  wire  decS_isNaR; // @[PositAdder.scala 52:32]
  wire  _T_886; // @[PositAdder.scala 53:33]
  wire  _T_887; // @[PositAdder.scala 53:21]
  wire  _T_888; // @[PositAdder.scala 53:52]
  wire  decS_isZero; // @[PositAdder.scala 53:37]
  wire [1:0] _T_890; // @[PositAdder.scala 54:33]
  wire  _T_891; // @[PositAdder.scala 54:49]
  wire  _T_892; // @[PositAdder.scala 54:63]
  wire  _T_893; // @[PositAdder.scala 54:53]
  wire [8:0] _GEN_6; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  wire [8:0] decS_scale; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  wire [2:0] _T_896; // @[convert.scala 46:61]
  wire [2:0] _T_897; // @[convert.scala 46:52]
  wire [2:0] _T_899; // @[convert.scala 46:42]
  wire [5:0] _T_900; // @[convert.scala 48:34]
  wire  _T_901; // @[convert.scala 49:36]
  wire [5:0] _T_903; // @[convert.scala 50:36]
  wire [5:0] _T_904; // @[convert.scala 50:36]
  wire [5:0] _T_905; // @[convert.scala 50:28]
  wire  _T_906; // @[convert.scala 51:31]
  wire  _T_907; // @[convert.scala 52:43]
  wire [29:0] _T_911; // @[Cat.scala 29:58]
  wire [5:0] _T_912; // @[Shift.scala 39:17]
  wire  _T_913; // @[Shift.scala 39:24]
  wire [4:0] _T_914; // @[Shift.scala 40:44]
  wire [13:0] _T_915; // @[Shift.scala 90:30]
  wire [15:0] _T_916; // @[Shift.scala 90:48]
  wire  _T_917; // @[Shift.scala 90:57]
  wire [13:0] _GEN_7; // @[Shift.scala 90:39]
  wire [13:0] _T_918; // @[Shift.scala 90:39]
  wire  _T_919; // @[Shift.scala 12:21]
  wire  _T_920; // @[Shift.scala 12:21]
  wire [15:0] _T_922; // @[Bitwise.scala 71:12]
  wire [29:0] _T_923; // @[Cat.scala 29:58]
  wire [29:0] _T_924; // @[Shift.scala 91:22]
  wire [3:0] _T_925; // @[Shift.scala 92:77]
  wire [21:0] _T_926; // @[Shift.scala 90:30]
  wire [7:0] _T_927; // @[Shift.scala 90:48]
  wire  _T_928; // @[Shift.scala 90:57]
  wire [21:0] _GEN_8; // @[Shift.scala 90:39]
  wire [21:0] _T_929; // @[Shift.scala 90:39]
  wire  _T_930; // @[Shift.scala 12:21]
  wire  _T_931; // @[Shift.scala 12:21]
  wire [7:0] _T_933; // @[Bitwise.scala 71:12]
  wire [29:0] _T_934; // @[Cat.scala 29:58]
  wire [29:0] _T_935; // @[Shift.scala 91:22]
  wire [2:0] _T_936; // @[Shift.scala 92:77]
  wire [25:0] _T_937; // @[Shift.scala 90:30]
  wire [3:0] _T_938; // @[Shift.scala 90:48]
  wire  _T_939; // @[Shift.scala 90:57]
  wire [25:0] _GEN_9; // @[Shift.scala 90:39]
  wire [25:0] _T_940; // @[Shift.scala 90:39]
  wire  _T_941; // @[Shift.scala 12:21]
  wire  _T_942; // @[Shift.scala 12:21]
  wire [3:0] _T_944; // @[Bitwise.scala 71:12]
  wire [29:0] _T_945; // @[Cat.scala 29:58]
  wire [29:0] _T_946; // @[Shift.scala 91:22]
  wire [1:0] _T_947; // @[Shift.scala 92:77]
  wire [27:0] _T_948; // @[Shift.scala 90:30]
  wire [1:0] _T_949; // @[Shift.scala 90:48]
  wire  _T_950; // @[Shift.scala 90:57]
  wire [27:0] _GEN_10; // @[Shift.scala 90:39]
  wire [27:0] _T_951; // @[Shift.scala 90:39]
  wire  _T_952; // @[Shift.scala 12:21]
  wire  _T_953; // @[Shift.scala 12:21]
  wire [1:0] _T_955; // @[Bitwise.scala 71:12]
  wire [29:0] _T_956; // @[Cat.scala 29:58]
  wire [29:0] _T_957; // @[Shift.scala 91:22]
  wire  _T_958; // @[Shift.scala 92:77]
  wire [28:0] _T_959; // @[Shift.scala 90:30]
  wire  _T_960; // @[Shift.scala 90:48]
  wire [28:0] _GEN_11; // @[Shift.scala 90:39]
  wire [28:0] _T_962; // @[Shift.scala 90:39]
  wire  _T_964; // @[Shift.scala 12:21]
  wire [29:0] _T_965; // @[Cat.scala 29:58]
  wire [29:0] _T_966; // @[Shift.scala 91:22]
  wire [29:0] _T_969; // @[Bitwise.scala 71:12]
  wire [29:0] _T_970; // @[Shift.scala 39:10]
  wire  _T_971; // @[convert.scala 55:31]
  wire  _T_972; // @[convert.scala 56:31]
  wire  _T_973; // @[convert.scala 57:31]
  wire  _T_974; // @[convert.scala 58:31]
  wire [26:0] _T_975; // @[convert.scala 59:69]
  wire  _T_976; // @[convert.scala 59:81]
  wire  _T_977; // @[convert.scala 59:50]
  wire  _T_979; // @[convert.scala 60:81]
  wire  _T_980; // @[convert.scala 61:44]
  wire  _T_981; // @[convert.scala 61:52]
  wire  _T_982; // @[convert.scala 61:36]
  wire  _T_983; // @[convert.scala 62:63]
  wire  _T_984; // @[convert.scala 62:103]
  wire  _T_985; // @[convert.scala 62:60]
  wire [26:0] _GEN_12; // @[convert.scala 63:56]
  wire [26:0] _T_988; // @[convert.scala 63:56]
  wire [27:0] _T_989; // @[Cat.scala 29:58]
  wire [27:0] _T_991; // @[Mux.scala 87:16]
  assign _T_1 = io_A[27]; // @[convert.scala 18:24]
  assign _T_2 = io_A[26]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[26:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[25:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[25:10]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[15:8]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[7:4]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9[3:2]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10 != 2'h0; // @[LZD.scala 39:14]
  assign _T_12 = _T_10[1]; // @[LZD.scala 39:21]
  assign _T_13 = _T_10[0]; // @[LZD.scala 39:30]
  assign _T_14 = ~ _T_13; // @[LZD.scala 39:27]
  assign _T_15 = _T_12 | _T_14; // @[LZD.scala 39:25]
  assign _T_16 = {_T_11,_T_15}; // @[Cat.scala 29:58]
  assign _T_17 = _T_9[1:0]; // @[LZD.scala 44:32]
  assign _T_18 = _T_17 != 2'h0; // @[LZD.scala 39:14]
  assign _T_19 = _T_17[1]; // @[LZD.scala 39:21]
  assign _T_20 = _T_17[0]; // @[LZD.scala 39:30]
  assign _T_21 = ~ _T_20; // @[LZD.scala 39:27]
  assign _T_22 = _T_19 | _T_21; // @[LZD.scala 39:25]
  assign _T_23 = {_T_18,_T_22}; // @[Cat.scala 29:58]
  assign _T_24 = _T_16[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23[1]; // @[Shift.scala 12:21]
  assign _T_26 = _T_24 | _T_25; // @[LZD.scala 49:16]
  assign _T_27 = ~ _T_25; // @[LZD.scala 49:27]
  assign _T_28 = _T_24 | _T_27; // @[LZD.scala 49:25]
  assign _T_29 = _T_16[0:0]; // @[LZD.scala 49:47]
  assign _T_30 = _T_23[0:0]; // @[LZD.scala 49:59]
  assign _T_31 = _T_24 ? _T_29 : _T_30; // @[LZD.scala 49:35]
  assign _T_33 = {_T_26,_T_28,_T_31}; // @[Cat.scala 29:58]
  assign _T_34 = _T_8[3:0]; // @[LZD.scala 44:32]
  assign _T_35 = _T_34[3:2]; // @[LZD.scala 43:32]
  assign _T_36 = _T_35 != 2'h0; // @[LZD.scala 39:14]
  assign _T_37 = _T_35[1]; // @[LZD.scala 39:21]
  assign _T_38 = _T_35[0]; // @[LZD.scala 39:30]
  assign _T_39 = ~ _T_38; // @[LZD.scala 39:27]
  assign _T_40 = _T_37 | _T_39; // @[LZD.scala 39:25]
  assign _T_41 = {_T_36,_T_40}; // @[Cat.scala 29:58]
  assign _T_42 = _T_34[1:0]; // @[LZD.scala 44:32]
  assign _T_43 = _T_42 != 2'h0; // @[LZD.scala 39:14]
  assign _T_44 = _T_42[1]; // @[LZD.scala 39:21]
  assign _T_45 = _T_42[0]; // @[LZD.scala 39:30]
  assign _T_46 = ~ _T_45; // @[LZD.scala 39:27]
  assign _T_47 = _T_44 | _T_46; // @[LZD.scala 39:25]
  assign _T_48 = {_T_43,_T_47}; // @[Cat.scala 29:58]
  assign _T_49 = _T_41[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48[1]; // @[Shift.scala 12:21]
  assign _T_51 = _T_49 | _T_50; // @[LZD.scala 49:16]
  assign _T_52 = ~ _T_50; // @[LZD.scala 49:27]
  assign _T_53 = _T_49 | _T_52; // @[LZD.scala 49:25]
  assign _T_54 = _T_41[0:0]; // @[LZD.scala 49:47]
  assign _T_55 = _T_48[0:0]; // @[LZD.scala 49:59]
  assign _T_56 = _T_49 ? _T_54 : _T_55; // @[LZD.scala 49:35]
  assign _T_58 = {_T_51,_T_53,_T_56}; // @[Cat.scala 29:58]
  assign _T_59 = _T_33[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58[2]; // @[Shift.scala 12:21]
  assign _T_61 = _T_59 | _T_60; // @[LZD.scala 49:16]
  assign _T_62 = ~ _T_60; // @[LZD.scala 49:27]
  assign _T_63 = _T_59 | _T_62; // @[LZD.scala 49:25]
  assign _T_64 = _T_33[1:0]; // @[LZD.scala 49:47]
  assign _T_65 = _T_58[1:0]; // @[LZD.scala 49:59]
  assign _T_66 = _T_59 ? _T_64 : _T_65; // @[LZD.scala 49:35]
  assign _T_68 = {_T_61,_T_63,_T_66}; // @[Cat.scala 29:58]
  assign _T_69 = _T_7[7:0]; // @[LZD.scala 44:32]
  assign _T_70 = _T_69[7:4]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70[3:2]; // @[LZD.scala 43:32]
  assign _T_72 = _T_71 != 2'h0; // @[LZD.scala 39:14]
  assign _T_73 = _T_71[1]; // @[LZD.scala 39:21]
  assign _T_74 = _T_71[0]; // @[LZD.scala 39:30]
  assign _T_75 = ~ _T_74; // @[LZD.scala 39:27]
  assign _T_76 = _T_73 | _T_75; // @[LZD.scala 39:25]
  assign _T_77 = {_T_72,_T_76}; // @[Cat.scala 29:58]
  assign _T_78 = _T_70[1:0]; // @[LZD.scala 44:32]
  assign _T_79 = _T_78 != 2'h0; // @[LZD.scala 39:14]
  assign _T_80 = _T_78[1]; // @[LZD.scala 39:21]
  assign _T_81 = _T_78[0]; // @[LZD.scala 39:30]
  assign _T_82 = ~ _T_81; // @[LZD.scala 39:27]
  assign _T_83 = _T_80 | _T_82; // @[LZD.scala 39:25]
  assign _T_84 = {_T_79,_T_83}; // @[Cat.scala 29:58]
  assign _T_85 = _T_77[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84[1]; // @[Shift.scala 12:21]
  assign _T_87 = _T_85 | _T_86; // @[LZD.scala 49:16]
  assign _T_88 = ~ _T_86; // @[LZD.scala 49:27]
  assign _T_89 = _T_85 | _T_88; // @[LZD.scala 49:25]
  assign _T_90 = _T_77[0:0]; // @[LZD.scala 49:47]
  assign _T_91 = _T_84[0:0]; // @[LZD.scala 49:59]
  assign _T_92 = _T_85 ? _T_90 : _T_91; // @[LZD.scala 49:35]
  assign _T_94 = {_T_87,_T_89,_T_92}; // @[Cat.scala 29:58]
  assign _T_95 = _T_69[3:0]; // @[LZD.scala 44:32]
  assign _T_96 = _T_95[3:2]; // @[LZD.scala 43:32]
  assign _T_97 = _T_96 != 2'h0; // @[LZD.scala 39:14]
  assign _T_98 = _T_96[1]; // @[LZD.scala 39:21]
  assign _T_99 = _T_96[0]; // @[LZD.scala 39:30]
  assign _T_100 = ~ _T_99; // @[LZD.scala 39:27]
  assign _T_101 = _T_98 | _T_100; // @[LZD.scala 39:25]
  assign _T_102 = {_T_97,_T_101}; // @[Cat.scala 29:58]
  assign _T_103 = _T_95[1:0]; // @[LZD.scala 44:32]
  assign _T_104 = _T_103 != 2'h0; // @[LZD.scala 39:14]
  assign _T_105 = _T_103[1]; // @[LZD.scala 39:21]
  assign _T_106 = _T_103[0]; // @[LZD.scala 39:30]
  assign _T_107 = ~ _T_106; // @[LZD.scala 39:27]
  assign _T_108 = _T_105 | _T_107; // @[LZD.scala 39:25]
  assign _T_109 = {_T_104,_T_108}; // @[Cat.scala 29:58]
  assign _T_110 = _T_102[1]; // @[Shift.scala 12:21]
  assign _T_111 = _T_109[1]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110 | _T_111; // @[LZD.scala 49:16]
  assign _T_113 = ~ _T_111; // @[LZD.scala 49:27]
  assign _T_114 = _T_110 | _T_113; // @[LZD.scala 49:25]
  assign _T_115 = _T_102[0:0]; // @[LZD.scala 49:47]
  assign _T_116 = _T_109[0:0]; // @[LZD.scala 49:59]
  assign _T_117 = _T_110 ? _T_115 : _T_116; // @[LZD.scala 49:35]
  assign _T_119 = {_T_112,_T_114,_T_117}; // @[Cat.scala 29:58]
  assign _T_120 = _T_94[2]; // @[Shift.scala 12:21]
  assign _T_121 = _T_119[2]; // @[Shift.scala 12:21]
  assign _T_122 = _T_120 | _T_121; // @[LZD.scala 49:16]
  assign _T_123 = ~ _T_121; // @[LZD.scala 49:27]
  assign _T_124 = _T_120 | _T_123; // @[LZD.scala 49:25]
  assign _T_125 = _T_94[1:0]; // @[LZD.scala 49:47]
  assign _T_126 = _T_119[1:0]; // @[LZD.scala 49:59]
  assign _T_127 = _T_120 ? _T_125 : _T_126; // @[LZD.scala 49:35]
  assign _T_129 = {_T_122,_T_124,_T_127}; // @[Cat.scala 29:58]
  assign _T_130 = _T_68[3]; // @[Shift.scala 12:21]
  assign _T_131 = _T_129[3]; // @[Shift.scala 12:21]
  assign _T_132 = _T_130 | _T_131; // @[LZD.scala 49:16]
  assign _T_133 = ~ _T_131; // @[LZD.scala 49:27]
  assign _T_134 = _T_130 | _T_133; // @[LZD.scala 49:25]
  assign _T_135 = _T_68[2:0]; // @[LZD.scala 49:47]
  assign _T_136 = _T_129[2:0]; // @[LZD.scala 49:59]
  assign _T_137 = _T_130 ? _T_135 : _T_136; // @[LZD.scala 49:35]
  assign _T_139 = {_T_132,_T_134,_T_137}; // @[Cat.scala 29:58]
  assign _T_140 = _T_6[9:0]; // @[LZD.scala 44:32]
  assign _T_141 = _T_140[9:2]; // @[LZD.scala 43:32]
  assign _T_142 = _T_141[7:4]; // @[LZD.scala 43:32]
  assign _T_143 = _T_142[3:2]; // @[LZD.scala 43:32]
  assign _T_144 = _T_143 != 2'h0; // @[LZD.scala 39:14]
  assign _T_145 = _T_143[1]; // @[LZD.scala 39:21]
  assign _T_146 = _T_143[0]; // @[LZD.scala 39:30]
  assign _T_147 = ~ _T_146; // @[LZD.scala 39:27]
  assign _T_148 = _T_145 | _T_147; // @[LZD.scala 39:25]
  assign _T_149 = {_T_144,_T_148}; // @[Cat.scala 29:58]
  assign _T_150 = _T_142[1:0]; // @[LZD.scala 44:32]
  assign _T_151 = _T_150 != 2'h0; // @[LZD.scala 39:14]
  assign _T_152 = _T_150[1]; // @[LZD.scala 39:21]
  assign _T_153 = _T_150[0]; // @[LZD.scala 39:30]
  assign _T_154 = ~ _T_153; // @[LZD.scala 39:27]
  assign _T_155 = _T_152 | _T_154; // @[LZD.scala 39:25]
  assign _T_156 = {_T_151,_T_155}; // @[Cat.scala 29:58]
  assign _T_157 = _T_149[1]; // @[Shift.scala 12:21]
  assign _T_158 = _T_156[1]; // @[Shift.scala 12:21]
  assign _T_159 = _T_157 | _T_158; // @[LZD.scala 49:16]
  assign _T_160 = ~ _T_158; // @[LZD.scala 49:27]
  assign _T_161 = _T_157 | _T_160; // @[LZD.scala 49:25]
  assign _T_162 = _T_149[0:0]; // @[LZD.scala 49:47]
  assign _T_163 = _T_156[0:0]; // @[LZD.scala 49:59]
  assign _T_164 = _T_157 ? _T_162 : _T_163; // @[LZD.scala 49:35]
  assign _T_166 = {_T_159,_T_161,_T_164}; // @[Cat.scala 29:58]
  assign _T_167 = _T_141[3:0]; // @[LZD.scala 44:32]
  assign _T_168 = _T_167[3:2]; // @[LZD.scala 43:32]
  assign _T_169 = _T_168 != 2'h0; // @[LZD.scala 39:14]
  assign _T_170 = _T_168[1]; // @[LZD.scala 39:21]
  assign _T_171 = _T_168[0]; // @[LZD.scala 39:30]
  assign _T_172 = ~ _T_171; // @[LZD.scala 39:27]
  assign _T_173 = _T_170 | _T_172; // @[LZD.scala 39:25]
  assign _T_174 = {_T_169,_T_173}; // @[Cat.scala 29:58]
  assign _T_175 = _T_167[1:0]; // @[LZD.scala 44:32]
  assign _T_176 = _T_175 != 2'h0; // @[LZD.scala 39:14]
  assign _T_177 = _T_175[1]; // @[LZD.scala 39:21]
  assign _T_178 = _T_175[0]; // @[LZD.scala 39:30]
  assign _T_179 = ~ _T_178; // @[LZD.scala 39:27]
  assign _T_180 = _T_177 | _T_179; // @[LZD.scala 39:25]
  assign _T_181 = {_T_176,_T_180}; // @[Cat.scala 29:58]
  assign _T_182 = _T_174[1]; // @[Shift.scala 12:21]
  assign _T_183 = _T_181[1]; // @[Shift.scala 12:21]
  assign _T_184 = _T_182 | _T_183; // @[LZD.scala 49:16]
  assign _T_185 = ~ _T_183; // @[LZD.scala 49:27]
  assign _T_186 = _T_182 | _T_185; // @[LZD.scala 49:25]
  assign _T_187 = _T_174[0:0]; // @[LZD.scala 49:47]
  assign _T_188 = _T_181[0:0]; // @[LZD.scala 49:59]
  assign _T_189 = _T_182 ? _T_187 : _T_188; // @[LZD.scala 49:35]
  assign _T_191 = {_T_184,_T_186,_T_189}; // @[Cat.scala 29:58]
  assign _T_192 = _T_166[2]; // @[Shift.scala 12:21]
  assign _T_193 = _T_191[2]; // @[Shift.scala 12:21]
  assign _T_194 = _T_192 | _T_193; // @[LZD.scala 49:16]
  assign _T_195 = ~ _T_193; // @[LZD.scala 49:27]
  assign _T_196 = _T_192 | _T_195; // @[LZD.scala 49:25]
  assign _T_197 = _T_166[1:0]; // @[LZD.scala 49:47]
  assign _T_198 = _T_191[1:0]; // @[LZD.scala 49:59]
  assign _T_199 = _T_192 ? _T_197 : _T_198; // @[LZD.scala 49:35]
  assign _T_201 = {_T_194,_T_196,_T_199}; // @[Cat.scala 29:58]
  assign _T_202 = _T_140[1:0]; // @[LZD.scala 44:32]
  assign _T_203 = _T_202 != 2'h0; // @[LZD.scala 39:14]
  assign _T_204 = _T_202[1]; // @[LZD.scala 39:21]
  assign _T_205 = _T_202[0]; // @[LZD.scala 39:30]
  assign _T_206 = ~ _T_205; // @[LZD.scala 39:27]
  assign _T_207 = _T_204 | _T_206; // @[LZD.scala 39:25]
  assign _T_209 = _T_201[3]; // @[Shift.scala 12:21]
  assign _T_211 = {1'h1,_T_203,_T_207}; // @[Cat.scala 29:58]
  assign _T_212 = _T_201[2:0]; // @[LZD.scala 55:32]
  assign _T_213 = _T_209 ? _T_212 : _T_211; // @[LZD.scala 55:20]
  assign _T_214 = {_T_209,_T_213}; // @[Cat.scala 29:58]
  assign _T_215 = _T_139[4]; // @[Shift.scala 12:21]
  assign _T_217 = _T_139[3:0]; // @[LZD.scala 55:32]
  assign _T_218 = _T_215 ? _T_217 : _T_214; // @[LZD.scala 55:20]
  assign _T_219 = {_T_215,_T_218}; // @[Cat.scala 29:58]
  assign _T_220 = ~ _T_219; // @[convert.scala 21:22]
  assign _T_221 = io_A[24:0]; // @[convert.scala 22:36]
  assign _T_222 = _T_220 < 5'h19; // @[Shift.scala 16:24]
  assign _T_224 = _T_220[4]; // @[Shift.scala 12:21]
  assign _T_225 = _T_221[8:0]; // @[Shift.scala 64:52]
  assign _T_227 = {_T_225,16'h0}; // @[Cat.scala 29:58]
  assign _T_228 = _T_224 ? _T_227 : _T_221; // @[Shift.scala 64:27]
  assign _T_229 = _T_220[3:0]; // @[Shift.scala 66:70]
  assign _T_230 = _T_229[3]; // @[Shift.scala 12:21]
  assign _T_231 = _T_228[16:0]; // @[Shift.scala 64:52]
  assign _T_233 = {_T_231,8'h0}; // @[Cat.scala 29:58]
  assign _T_234 = _T_230 ? _T_233 : _T_228; // @[Shift.scala 64:27]
  assign _T_235 = _T_229[2:0]; // @[Shift.scala 66:70]
  assign _T_236 = _T_235[2]; // @[Shift.scala 12:21]
  assign _T_237 = _T_234[20:0]; // @[Shift.scala 64:52]
  assign _T_239 = {_T_237,4'h0}; // @[Cat.scala 29:58]
  assign _T_240 = _T_236 ? _T_239 : _T_234; // @[Shift.scala 64:27]
  assign _T_241 = _T_235[1:0]; // @[Shift.scala 66:70]
  assign _T_242 = _T_241[1]; // @[Shift.scala 12:21]
  assign _T_243 = _T_240[22:0]; // @[Shift.scala 64:52]
  assign _T_245 = {_T_243,2'h0}; // @[Cat.scala 29:58]
  assign _T_246 = _T_242 ? _T_245 : _T_240; // @[Shift.scala 64:27]
  assign _T_247 = _T_241[0:0]; // @[Shift.scala 66:70]
  assign _T_249 = _T_246[23:0]; // @[Shift.scala 64:52]
  assign _T_250 = {_T_249,1'h0}; // @[Cat.scala 29:58]
  assign _T_251 = _T_247 ? _T_250 : _T_246; // @[Shift.scala 64:27]
  assign _T_252 = _T_222 ? _T_251 : 25'h0; // @[Shift.scala 16:10]
  assign _T_253 = _T_252[24:22]; // @[convert.scala 23:34]
  assign decA_fraction = _T_252[21:0]; // @[convert.scala 24:34]
  assign _T_255 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_257 = _T_3 ? _T_220 : _T_219; // @[convert.scala 25:42]
  assign _T_260 = ~ _T_253; // @[convert.scala 26:67]
  assign _T_261 = _T_1 ? _T_260 : _T_253; // @[convert.scala 26:51]
  assign _T_262 = {_T_255,_T_257,_T_261}; // @[Cat.scala 29:58]
  assign _T_264 = io_A[26:0]; // @[convert.scala 29:56]
  assign _T_265 = _T_264 != 27'h0; // @[convert.scala 29:60]
  assign _T_266 = ~ _T_265; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_266; // @[convert.scala 29:39]
  assign _T_269 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_269 & _T_266; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_262); // @[convert.scala 32:24]
  assign _T_278 = io_B[27]; // @[convert.scala 18:24]
  assign _T_279 = io_B[26]; // @[convert.scala 18:40]
  assign _T_280 = _T_278 ^ _T_279; // @[convert.scala 18:36]
  assign _T_281 = io_B[26:1]; // @[convert.scala 19:24]
  assign _T_282 = io_B[25:0]; // @[convert.scala 19:43]
  assign _T_283 = _T_281 ^ _T_282; // @[convert.scala 19:39]
  assign _T_284 = _T_283[25:10]; // @[LZD.scala 43:32]
  assign _T_285 = _T_284[15:8]; // @[LZD.scala 43:32]
  assign _T_286 = _T_285[7:4]; // @[LZD.scala 43:32]
  assign _T_287 = _T_286[3:2]; // @[LZD.scala 43:32]
  assign _T_288 = _T_287 != 2'h0; // @[LZD.scala 39:14]
  assign _T_289 = _T_287[1]; // @[LZD.scala 39:21]
  assign _T_290 = _T_287[0]; // @[LZD.scala 39:30]
  assign _T_291 = ~ _T_290; // @[LZD.scala 39:27]
  assign _T_292 = _T_289 | _T_291; // @[LZD.scala 39:25]
  assign _T_293 = {_T_288,_T_292}; // @[Cat.scala 29:58]
  assign _T_294 = _T_286[1:0]; // @[LZD.scala 44:32]
  assign _T_295 = _T_294 != 2'h0; // @[LZD.scala 39:14]
  assign _T_296 = _T_294[1]; // @[LZD.scala 39:21]
  assign _T_297 = _T_294[0]; // @[LZD.scala 39:30]
  assign _T_298 = ~ _T_297; // @[LZD.scala 39:27]
  assign _T_299 = _T_296 | _T_298; // @[LZD.scala 39:25]
  assign _T_300 = {_T_295,_T_299}; // @[Cat.scala 29:58]
  assign _T_301 = _T_293[1]; // @[Shift.scala 12:21]
  assign _T_302 = _T_300[1]; // @[Shift.scala 12:21]
  assign _T_303 = _T_301 | _T_302; // @[LZD.scala 49:16]
  assign _T_304 = ~ _T_302; // @[LZD.scala 49:27]
  assign _T_305 = _T_301 | _T_304; // @[LZD.scala 49:25]
  assign _T_306 = _T_293[0:0]; // @[LZD.scala 49:47]
  assign _T_307 = _T_300[0:0]; // @[LZD.scala 49:59]
  assign _T_308 = _T_301 ? _T_306 : _T_307; // @[LZD.scala 49:35]
  assign _T_310 = {_T_303,_T_305,_T_308}; // @[Cat.scala 29:58]
  assign _T_311 = _T_285[3:0]; // @[LZD.scala 44:32]
  assign _T_312 = _T_311[3:2]; // @[LZD.scala 43:32]
  assign _T_313 = _T_312 != 2'h0; // @[LZD.scala 39:14]
  assign _T_314 = _T_312[1]; // @[LZD.scala 39:21]
  assign _T_315 = _T_312[0]; // @[LZD.scala 39:30]
  assign _T_316 = ~ _T_315; // @[LZD.scala 39:27]
  assign _T_317 = _T_314 | _T_316; // @[LZD.scala 39:25]
  assign _T_318 = {_T_313,_T_317}; // @[Cat.scala 29:58]
  assign _T_319 = _T_311[1:0]; // @[LZD.scala 44:32]
  assign _T_320 = _T_319 != 2'h0; // @[LZD.scala 39:14]
  assign _T_321 = _T_319[1]; // @[LZD.scala 39:21]
  assign _T_322 = _T_319[0]; // @[LZD.scala 39:30]
  assign _T_323 = ~ _T_322; // @[LZD.scala 39:27]
  assign _T_324 = _T_321 | _T_323; // @[LZD.scala 39:25]
  assign _T_325 = {_T_320,_T_324}; // @[Cat.scala 29:58]
  assign _T_326 = _T_318[1]; // @[Shift.scala 12:21]
  assign _T_327 = _T_325[1]; // @[Shift.scala 12:21]
  assign _T_328 = _T_326 | _T_327; // @[LZD.scala 49:16]
  assign _T_329 = ~ _T_327; // @[LZD.scala 49:27]
  assign _T_330 = _T_326 | _T_329; // @[LZD.scala 49:25]
  assign _T_331 = _T_318[0:0]; // @[LZD.scala 49:47]
  assign _T_332 = _T_325[0:0]; // @[LZD.scala 49:59]
  assign _T_333 = _T_326 ? _T_331 : _T_332; // @[LZD.scala 49:35]
  assign _T_335 = {_T_328,_T_330,_T_333}; // @[Cat.scala 29:58]
  assign _T_336 = _T_310[2]; // @[Shift.scala 12:21]
  assign _T_337 = _T_335[2]; // @[Shift.scala 12:21]
  assign _T_338 = _T_336 | _T_337; // @[LZD.scala 49:16]
  assign _T_339 = ~ _T_337; // @[LZD.scala 49:27]
  assign _T_340 = _T_336 | _T_339; // @[LZD.scala 49:25]
  assign _T_341 = _T_310[1:0]; // @[LZD.scala 49:47]
  assign _T_342 = _T_335[1:0]; // @[LZD.scala 49:59]
  assign _T_343 = _T_336 ? _T_341 : _T_342; // @[LZD.scala 49:35]
  assign _T_345 = {_T_338,_T_340,_T_343}; // @[Cat.scala 29:58]
  assign _T_346 = _T_284[7:0]; // @[LZD.scala 44:32]
  assign _T_347 = _T_346[7:4]; // @[LZD.scala 43:32]
  assign _T_348 = _T_347[3:2]; // @[LZD.scala 43:32]
  assign _T_349 = _T_348 != 2'h0; // @[LZD.scala 39:14]
  assign _T_350 = _T_348[1]; // @[LZD.scala 39:21]
  assign _T_351 = _T_348[0]; // @[LZD.scala 39:30]
  assign _T_352 = ~ _T_351; // @[LZD.scala 39:27]
  assign _T_353 = _T_350 | _T_352; // @[LZD.scala 39:25]
  assign _T_354 = {_T_349,_T_353}; // @[Cat.scala 29:58]
  assign _T_355 = _T_347[1:0]; // @[LZD.scala 44:32]
  assign _T_356 = _T_355 != 2'h0; // @[LZD.scala 39:14]
  assign _T_357 = _T_355[1]; // @[LZD.scala 39:21]
  assign _T_358 = _T_355[0]; // @[LZD.scala 39:30]
  assign _T_359 = ~ _T_358; // @[LZD.scala 39:27]
  assign _T_360 = _T_357 | _T_359; // @[LZD.scala 39:25]
  assign _T_361 = {_T_356,_T_360}; // @[Cat.scala 29:58]
  assign _T_362 = _T_354[1]; // @[Shift.scala 12:21]
  assign _T_363 = _T_361[1]; // @[Shift.scala 12:21]
  assign _T_364 = _T_362 | _T_363; // @[LZD.scala 49:16]
  assign _T_365 = ~ _T_363; // @[LZD.scala 49:27]
  assign _T_366 = _T_362 | _T_365; // @[LZD.scala 49:25]
  assign _T_367 = _T_354[0:0]; // @[LZD.scala 49:47]
  assign _T_368 = _T_361[0:0]; // @[LZD.scala 49:59]
  assign _T_369 = _T_362 ? _T_367 : _T_368; // @[LZD.scala 49:35]
  assign _T_371 = {_T_364,_T_366,_T_369}; // @[Cat.scala 29:58]
  assign _T_372 = _T_346[3:0]; // @[LZD.scala 44:32]
  assign _T_373 = _T_372[3:2]; // @[LZD.scala 43:32]
  assign _T_374 = _T_373 != 2'h0; // @[LZD.scala 39:14]
  assign _T_375 = _T_373[1]; // @[LZD.scala 39:21]
  assign _T_376 = _T_373[0]; // @[LZD.scala 39:30]
  assign _T_377 = ~ _T_376; // @[LZD.scala 39:27]
  assign _T_378 = _T_375 | _T_377; // @[LZD.scala 39:25]
  assign _T_379 = {_T_374,_T_378}; // @[Cat.scala 29:58]
  assign _T_380 = _T_372[1:0]; // @[LZD.scala 44:32]
  assign _T_381 = _T_380 != 2'h0; // @[LZD.scala 39:14]
  assign _T_382 = _T_380[1]; // @[LZD.scala 39:21]
  assign _T_383 = _T_380[0]; // @[LZD.scala 39:30]
  assign _T_384 = ~ _T_383; // @[LZD.scala 39:27]
  assign _T_385 = _T_382 | _T_384; // @[LZD.scala 39:25]
  assign _T_386 = {_T_381,_T_385}; // @[Cat.scala 29:58]
  assign _T_387 = _T_379[1]; // @[Shift.scala 12:21]
  assign _T_388 = _T_386[1]; // @[Shift.scala 12:21]
  assign _T_389 = _T_387 | _T_388; // @[LZD.scala 49:16]
  assign _T_390 = ~ _T_388; // @[LZD.scala 49:27]
  assign _T_391 = _T_387 | _T_390; // @[LZD.scala 49:25]
  assign _T_392 = _T_379[0:0]; // @[LZD.scala 49:47]
  assign _T_393 = _T_386[0:0]; // @[LZD.scala 49:59]
  assign _T_394 = _T_387 ? _T_392 : _T_393; // @[LZD.scala 49:35]
  assign _T_396 = {_T_389,_T_391,_T_394}; // @[Cat.scala 29:58]
  assign _T_397 = _T_371[2]; // @[Shift.scala 12:21]
  assign _T_398 = _T_396[2]; // @[Shift.scala 12:21]
  assign _T_399 = _T_397 | _T_398; // @[LZD.scala 49:16]
  assign _T_400 = ~ _T_398; // @[LZD.scala 49:27]
  assign _T_401 = _T_397 | _T_400; // @[LZD.scala 49:25]
  assign _T_402 = _T_371[1:0]; // @[LZD.scala 49:47]
  assign _T_403 = _T_396[1:0]; // @[LZD.scala 49:59]
  assign _T_404 = _T_397 ? _T_402 : _T_403; // @[LZD.scala 49:35]
  assign _T_406 = {_T_399,_T_401,_T_404}; // @[Cat.scala 29:58]
  assign _T_407 = _T_345[3]; // @[Shift.scala 12:21]
  assign _T_408 = _T_406[3]; // @[Shift.scala 12:21]
  assign _T_409 = _T_407 | _T_408; // @[LZD.scala 49:16]
  assign _T_410 = ~ _T_408; // @[LZD.scala 49:27]
  assign _T_411 = _T_407 | _T_410; // @[LZD.scala 49:25]
  assign _T_412 = _T_345[2:0]; // @[LZD.scala 49:47]
  assign _T_413 = _T_406[2:0]; // @[LZD.scala 49:59]
  assign _T_414 = _T_407 ? _T_412 : _T_413; // @[LZD.scala 49:35]
  assign _T_416 = {_T_409,_T_411,_T_414}; // @[Cat.scala 29:58]
  assign _T_417 = _T_283[9:0]; // @[LZD.scala 44:32]
  assign _T_418 = _T_417[9:2]; // @[LZD.scala 43:32]
  assign _T_419 = _T_418[7:4]; // @[LZD.scala 43:32]
  assign _T_420 = _T_419[3:2]; // @[LZD.scala 43:32]
  assign _T_421 = _T_420 != 2'h0; // @[LZD.scala 39:14]
  assign _T_422 = _T_420[1]; // @[LZD.scala 39:21]
  assign _T_423 = _T_420[0]; // @[LZD.scala 39:30]
  assign _T_424 = ~ _T_423; // @[LZD.scala 39:27]
  assign _T_425 = _T_422 | _T_424; // @[LZD.scala 39:25]
  assign _T_426 = {_T_421,_T_425}; // @[Cat.scala 29:58]
  assign _T_427 = _T_419[1:0]; // @[LZD.scala 44:32]
  assign _T_428 = _T_427 != 2'h0; // @[LZD.scala 39:14]
  assign _T_429 = _T_427[1]; // @[LZD.scala 39:21]
  assign _T_430 = _T_427[0]; // @[LZD.scala 39:30]
  assign _T_431 = ~ _T_430; // @[LZD.scala 39:27]
  assign _T_432 = _T_429 | _T_431; // @[LZD.scala 39:25]
  assign _T_433 = {_T_428,_T_432}; // @[Cat.scala 29:58]
  assign _T_434 = _T_426[1]; // @[Shift.scala 12:21]
  assign _T_435 = _T_433[1]; // @[Shift.scala 12:21]
  assign _T_436 = _T_434 | _T_435; // @[LZD.scala 49:16]
  assign _T_437 = ~ _T_435; // @[LZD.scala 49:27]
  assign _T_438 = _T_434 | _T_437; // @[LZD.scala 49:25]
  assign _T_439 = _T_426[0:0]; // @[LZD.scala 49:47]
  assign _T_440 = _T_433[0:0]; // @[LZD.scala 49:59]
  assign _T_441 = _T_434 ? _T_439 : _T_440; // @[LZD.scala 49:35]
  assign _T_443 = {_T_436,_T_438,_T_441}; // @[Cat.scala 29:58]
  assign _T_444 = _T_418[3:0]; // @[LZD.scala 44:32]
  assign _T_445 = _T_444[3:2]; // @[LZD.scala 43:32]
  assign _T_446 = _T_445 != 2'h0; // @[LZD.scala 39:14]
  assign _T_447 = _T_445[1]; // @[LZD.scala 39:21]
  assign _T_448 = _T_445[0]; // @[LZD.scala 39:30]
  assign _T_449 = ~ _T_448; // @[LZD.scala 39:27]
  assign _T_450 = _T_447 | _T_449; // @[LZD.scala 39:25]
  assign _T_451 = {_T_446,_T_450}; // @[Cat.scala 29:58]
  assign _T_452 = _T_444[1:0]; // @[LZD.scala 44:32]
  assign _T_453 = _T_452 != 2'h0; // @[LZD.scala 39:14]
  assign _T_454 = _T_452[1]; // @[LZD.scala 39:21]
  assign _T_455 = _T_452[0]; // @[LZD.scala 39:30]
  assign _T_456 = ~ _T_455; // @[LZD.scala 39:27]
  assign _T_457 = _T_454 | _T_456; // @[LZD.scala 39:25]
  assign _T_458 = {_T_453,_T_457}; // @[Cat.scala 29:58]
  assign _T_459 = _T_451[1]; // @[Shift.scala 12:21]
  assign _T_460 = _T_458[1]; // @[Shift.scala 12:21]
  assign _T_461 = _T_459 | _T_460; // @[LZD.scala 49:16]
  assign _T_462 = ~ _T_460; // @[LZD.scala 49:27]
  assign _T_463 = _T_459 | _T_462; // @[LZD.scala 49:25]
  assign _T_464 = _T_451[0:0]; // @[LZD.scala 49:47]
  assign _T_465 = _T_458[0:0]; // @[LZD.scala 49:59]
  assign _T_466 = _T_459 ? _T_464 : _T_465; // @[LZD.scala 49:35]
  assign _T_468 = {_T_461,_T_463,_T_466}; // @[Cat.scala 29:58]
  assign _T_469 = _T_443[2]; // @[Shift.scala 12:21]
  assign _T_470 = _T_468[2]; // @[Shift.scala 12:21]
  assign _T_471 = _T_469 | _T_470; // @[LZD.scala 49:16]
  assign _T_472 = ~ _T_470; // @[LZD.scala 49:27]
  assign _T_473 = _T_469 | _T_472; // @[LZD.scala 49:25]
  assign _T_474 = _T_443[1:0]; // @[LZD.scala 49:47]
  assign _T_475 = _T_468[1:0]; // @[LZD.scala 49:59]
  assign _T_476 = _T_469 ? _T_474 : _T_475; // @[LZD.scala 49:35]
  assign _T_478 = {_T_471,_T_473,_T_476}; // @[Cat.scala 29:58]
  assign _T_479 = _T_417[1:0]; // @[LZD.scala 44:32]
  assign _T_480 = _T_479 != 2'h0; // @[LZD.scala 39:14]
  assign _T_481 = _T_479[1]; // @[LZD.scala 39:21]
  assign _T_482 = _T_479[0]; // @[LZD.scala 39:30]
  assign _T_483 = ~ _T_482; // @[LZD.scala 39:27]
  assign _T_484 = _T_481 | _T_483; // @[LZD.scala 39:25]
  assign _T_486 = _T_478[3]; // @[Shift.scala 12:21]
  assign _T_488 = {1'h1,_T_480,_T_484}; // @[Cat.scala 29:58]
  assign _T_489 = _T_478[2:0]; // @[LZD.scala 55:32]
  assign _T_490 = _T_486 ? _T_489 : _T_488; // @[LZD.scala 55:20]
  assign _T_491 = {_T_486,_T_490}; // @[Cat.scala 29:58]
  assign _T_492 = _T_416[4]; // @[Shift.scala 12:21]
  assign _T_494 = _T_416[3:0]; // @[LZD.scala 55:32]
  assign _T_495 = _T_492 ? _T_494 : _T_491; // @[LZD.scala 55:20]
  assign _T_496 = {_T_492,_T_495}; // @[Cat.scala 29:58]
  assign _T_497 = ~ _T_496; // @[convert.scala 21:22]
  assign _T_498 = io_B[24:0]; // @[convert.scala 22:36]
  assign _T_499 = _T_497 < 5'h19; // @[Shift.scala 16:24]
  assign _T_501 = _T_497[4]; // @[Shift.scala 12:21]
  assign _T_502 = _T_498[8:0]; // @[Shift.scala 64:52]
  assign _T_504 = {_T_502,16'h0}; // @[Cat.scala 29:58]
  assign _T_505 = _T_501 ? _T_504 : _T_498; // @[Shift.scala 64:27]
  assign _T_506 = _T_497[3:0]; // @[Shift.scala 66:70]
  assign _T_507 = _T_506[3]; // @[Shift.scala 12:21]
  assign _T_508 = _T_505[16:0]; // @[Shift.scala 64:52]
  assign _T_510 = {_T_508,8'h0}; // @[Cat.scala 29:58]
  assign _T_511 = _T_507 ? _T_510 : _T_505; // @[Shift.scala 64:27]
  assign _T_512 = _T_506[2:0]; // @[Shift.scala 66:70]
  assign _T_513 = _T_512[2]; // @[Shift.scala 12:21]
  assign _T_514 = _T_511[20:0]; // @[Shift.scala 64:52]
  assign _T_516 = {_T_514,4'h0}; // @[Cat.scala 29:58]
  assign _T_517 = _T_513 ? _T_516 : _T_511; // @[Shift.scala 64:27]
  assign _T_518 = _T_512[1:0]; // @[Shift.scala 66:70]
  assign _T_519 = _T_518[1]; // @[Shift.scala 12:21]
  assign _T_520 = _T_517[22:0]; // @[Shift.scala 64:52]
  assign _T_522 = {_T_520,2'h0}; // @[Cat.scala 29:58]
  assign _T_523 = _T_519 ? _T_522 : _T_517; // @[Shift.scala 64:27]
  assign _T_524 = _T_518[0:0]; // @[Shift.scala 66:70]
  assign _T_526 = _T_523[23:0]; // @[Shift.scala 64:52]
  assign _T_527 = {_T_526,1'h0}; // @[Cat.scala 29:58]
  assign _T_528 = _T_524 ? _T_527 : _T_523; // @[Shift.scala 64:27]
  assign _T_529 = _T_499 ? _T_528 : 25'h0; // @[Shift.scala 16:10]
  assign _T_530 = _T_529[24:22]; // @[convert.scala 23:34]
  assign decB_fraction = _T_529[21:0]; // @[convert.scala 24:34]
  assign _T_532 = _T_280 == 1'h0; // @[convert.scala 25:26]
  assign _T_534 = _T_280 ? _T_497 : _T_496; // @[convert.scala 25:42]
  assign _T_537 = ~ _T_530; // @[convert.scala 26:67]
  assign _T_538 = _T_278 ? _T_537 : _T_530; // @[convert.scala 26:51]
  assign _T_539 = {_T_532,_T_534,_T_538}; // @[Cat.scala 29:58]
  assign _T_541 = io_B[26:0]; // @[convert.scala 29:56]
  assign _T_542 = _T_541 != 27'h0; // @[convert.scala 29:60]
  assign _T_543 = ~ _T_542; // @[convert.scala 29:41]
  assign decB_isNaR = _T_278 & _T_543; // @[convert.scala 29:39]
  assign _T_546 = _T_278 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_546 & _T_543; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_539); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[PositAdder.scala 24:32]
  assign greaterSign = aGTb ? _T_1 : _T_278; // @[PositAdder.scala 25:24]
  assign smallerSign = aGTb ? _T_278 : _T_1; // @[PositAdder.scala 26:24]
  assign greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[PositAdder.scala 27:24]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[PositAdder.scala 28:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[PositAdder.scala 29:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[PositAdder.scala 30:24]
  assign _T_555 = $signed(greaterExp) - $signed(smallerExp); // @[PositAdder.scala 31:32]
  assign scale_diff = $signed(_T_555); // @[PositAdder.scala 31:32]
  assign _T_556 = ~ greaterSign; // @[PositAdder.scala 32:38]
  assign greaterSig = {greaterSign,_T_556,greaterFrac}; // @[Cat.scala 29:58]
  assign _T_558 = ~ smallerSign; // @[PositAdder.scala 33:38]
  assign _T_561 = {smallerSign,_T_558,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_562 = $unsigned(scale_diff); // @[PositAdder.scala 34:68]
  assign _T_563 = _T_562 < 9'h1b; // @[Shift.scala 39:24]
  assign _T_564 = _T_562[4:0]; // @[Shift.scala 40:44]
  assign _T_565 = _T_561[26:16]; // @[Shift.scala 90:30]
  assign _T_566 = _T_561[15:0]; // @[Shift.scala 90:48]
  assign _T_567 = _T_566 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{10'd0}, _T_567}; // @[Shift.scala 90:39]
  assign _T_568 = _T_565 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_569 = _T_564[4]; // @[Shift.scala 12:21]
  assign _T_570 = _T_561[26]; // @[Shift.scala 12:21]
  assign _T_572 = _T_570 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_573 = {_T_572,_T_568}; // @[Cat.scala 29:58]
  assign _T_574 = _T_569 ? _T_573 : _T_561; // @[Shift.scala 91:22]
  assign _T_575 = _T_564[3:0]; // @[Shift.scala 92:77]
  assign _T_576 = _T_574[26:8]; // @[Shift.scala 90:30]
  assign _T_577 = _T_574[7:0]; // @[Shift.scala 90:48]
  assign _T_578 = _T_577 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{18'd0}, _T_578}; // @[Shift.scala 90:39]
  assign _T_579 = _T_576 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_580 = _T_575[3]; // @[Shift.scala 12:21]
  assign _T_581 = _T_574[26]; // @[Shift.scala 12:21]
  assign _T_583 = _T_581 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_584 = {_T_583,_T_579}; // @[Cat.scala 29:58]
  assign _T_585 = _T_580 ? _T_584 : _T_574; // @[Shift.scala 91:22]
  assign _T_586 = _T_575[2:0]; // @[Shift.scala 92:77]
  assign _T_587 = _T_585[26:4]; // @[Shift.scala 90:30]
  assign _T_588 = _T_585[3:0]; // @[Shift.scala 90:48]
  assign _T_589 = _T_588 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{22'd0}, _T_589}; // @[Shift.scala 90:39]
  assign _T_590 = _T_587 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_591 = _T_586[2]; // @[Shift.scala 12:21]
  assign _T_592 = _T_585[26]; // @[Shift.scala 12:21]
  assign _T_594 = _T_592 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_595 = {_T_594,_T_590}; // @[Cat.scala 29:58]
  assign _T_596 = _T_591 ? _T_595 : _T_585; // @[Shift.scala 91:22]
  assign _T_597 = _T_586[1:0]; // @[Shift.scala 92:77]
  assign _T_598 = _T_596[26:2]; // @[Shift.scala 90:30]
  assign _T_599 = _T_596[1:0]; // @[Shift.scala 90:48]
  assign _T_600 = _T_599 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_3 = {{24'd0}, _T_600}; // @[Shift.scala 90:39]
  assign _T_601 = _T_598 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_602 = _T_597[1]; // @[Shift.scala 12:21]
  assign _T_603 = _T_596[26]; // @[Shift.scala 12:21]
  assign _T_605 = _T_603 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_606 = {_T_605,_T_601}; // @[Cat.scala 29:58]
  assign _T_607 = _T_602 ? _T_606 : _T_596; // @[Shift.scala 91:22]
  assign _T_608 = _T_597[0:0]; // @[Shift.scala 92:77]
  assign _T_609 = _T_607[26:1]; // @[Shift.scala 90:30]
  assign _T_610 = _T_607[0:0]; // @[Shift.scala 90:48]
  assign _GEN_4 = {{25'd0}, _T_610}; // @[Shift.scala 90:39]
  assign _T_612 = _T_609 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_614 = _T_607[26]; // @[Shift.scala 12:21]
  assign _T_615 = {_T_614,_T_612}; // @[Cat.scala 29:58]
  assign _T_616 = _T_608 ? _T_615 : _T_607; // @[Shift.scala 91:22]
  assign _T_619 = _T_570 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_563 ? _T_616 : _T_619; // @[Shift.scala 39:10]
  assign _T_620 = smallerSig[26:3]; // @[PositAdder.scala 35:45]
  assign rawSumSig = greaterSig + _T_620; // @[PositAdder.scala 35:32]
  assign _T_621 = _T_1 ^ _T_278; // @[PositAdder.scala 36:31]
  assign _T_622 = rawSumSig[24:24]; // @[PositAdder.scala 36:59]
  assign sumSign = _T_621 ^ _T_622; // @[PositAdder.scala 36:43]
  assign _T_623 = greaterSig + _T_620; // @[PositAdder.scala 37:48]
  assign _T_624 = smallerSig[2:0]; // @[PositAdder.scala 37:63]
  assign signSumSig = {sumSign,_T_623,_T_624}; // @[Cat.scala 29:58]
  assign _T_626 = signSumSig[27:1]; // @[PositAdder.scala 39:31]
  assign _T_627 = signSumSig[26:0]; // @[PositAdder.scala 39:66]
  assign sumXor = _T_626 ^ _T_627; // @[PositAdder.scala 39:49]
  assign _T_628 = sumXor[26:11]; // @[LZD.scala 43:32]
  assign _T_629 = _T_628[15:8]; // @[LZD.scala 43:32]
  assign _T_630 = _T_629[7:4]; // @[LZD.scala 43:32]
  assign _T_631 = _T_630[3:2]; // @[LZD.scala 43:32]
  assign _T_632 = _T_631 != 2'h0; // @[LZD.scala 39:14]
  assign _T_633 = _T_631[1]; // @[LZD.scala 39:21]
  assign _T_634 = _T_631[0]; // @[LZD.scala 39:30]
  assign _T_635 = ~ _T_634; // @[LZD.scala 39:27]
  assign _T_636 = _T_633 | _T_635; // @[LZD.scala 39:25]
  assign _T_637 = {_T_632,_T_636}; // @[Cat.scala 29:58]
  assign _T_638 = _T_630[1:0]; // @[LZD.scala 44:32]
  assign _T_639 = _T_638 != 2'h0; // @[LZD.scala 39:14]
  assign _T_640 = _T_638[1]; // @[LZD.scala 39:21]
  assign _T_641 = _T_638[0]; // @[LZD.scala 39:30]
  assign _T_642 = ~ _T_641; // @[LZD.scala 39:27]
  assign _T_643 = _T_640 | _T_642; // @[LZD.scala 39:25]
  assign _T_644 = {_T_639,_T_643}; // @[Cat.scala 29:58]
  assign _T_645 = _T_637[1]; // @[Shift.scala 12:21]
  assign _T_646 = _T_644[1]; // @[Shift.scala 12:21]
  assign _T_647 = _T_645 | _T_646; // @[LZD.scala 49:16]
  assign _T_648 = ~ _T_646; // @[LZD.scala 49:27]
  assign _T_649 = _T_645 | _T_648; // @[LZD.scala 49:25]
  assign _T_650 = _T_637[0:0]; // @[LZD.scala 49:47]
  assign _T_651 = _T_644[0:0]; // @[LZD.scala 49:59]
  assign _T_652 = _T_645 ? _T_650 : _T_651; // @[LZD.scala 49:35]
  assign _T_654 = {_T_647,_T_649,_T_652}; // @[Cat.scala 29:58]
  assign _T_655 = _T_629[3:0]; // @[LZD.scala 44:32]
  assign _T_656 = _T_655[3:2]; // @[LZD.scala 43:32]
  assign _T_657 = _T_656 != 2'h0; // @[LZD.scala 39:14]
  assign _T_658 = _T_656[1]; // @[LZD.scala 39:21]
  assign _T_659 = _T_656[0]; // @[LZD.scala 39:30]
  assign _T_660 = ~ _T_659; // @[LZD.scala 39:27]
  assign _T_661 = _T_658 | _T_660; // @[LZD.scala 39:25]
  assign _T_662 = {_T_657,_T_661}; // @[Cat.scala 29:58]
  assign _T_663 = _T_655[1:0]; // @[LZD.scala 44:32]
  assign _T_664 = _T_663 != 2'h0; // @[LZD.scala 39:14]
  assign _T_665 = _T_663[1]; // @[LZD.scala 39:21]
  assign _T_666 = _T_663[0]; // @[LZD.scala 39:30]
  assign _T_667 = ~ _T_666; // @[LZD.scala 39:27]
  assign _T_668 = _T_665 | _T_667; // @[LZD.scala 39:25]
  assign _T_669 = {_T_664,_T_668}; // @[Cat.scala 29:58]
  assign _T_670 = _T_662[1]; // @[Shift.scala 12:21]
  assign _T_671 = _T_669[1]; // @[Shift.scala 12:21]
  assign _T_672 = _T_670 | _T_671; // @[LZD.scala 49:16]
  assign _T_673 = ~ _T_671; // @[LZD.scala 49:27]
  assign _T_674 = _T_670 | _T_673; // @[LZD.scala 49:25]
  assign _T_675 = _T_662[0:0]; // @[LZD.scala 49:47]
  assign _T_676 = _T_669[0:0]; // @[LZD.scala 49:59]
  assign _T_677 = _T_670 ? _T_675 : _T_676; // @[LZD.scala 49:35]
  assign _T_679 = {_T_672,_T_674,_T_677}; // @[Cat.scala 29:58]
  assign _T_680 = _T_654[2]; // @[Shift.scala 12:21]
  assign _T_681 = _T_679[2]; // @[Shift.scala 12:21]
  assign _T_682 = _T_680 | _T_681; // @[LZD.scala 49:16]
  assign _T_683 = ~ _T_681; // @[LZD.scala 49:27]
  assign _T_684 = _T_680 | _T_683; // @[LZD.scala 49:25]
  assign _T_685 = _T_654[1:0]; // @[LZD.scala 49:47]
  assign _T_686 = _T_679[1:0]; // @[LZD.scala 49:59]
  assign _T_687 = _T_680 ? _T_685 : _T_686; // @[LZD.scala 49:35]
  assign _T_689 = {_T_682,_T_684,_T_687}; // @[Cat.scala 29:58]
  assign _T_690 = _T_628[7:0]; // @[LZD.scala 44:32]
  assign _T_691 = _T_690[7:4]; // @[LZD.scala 43:32]
  assign _T_692 = _T_691[3:2]; // @[LZD.scala 43:32]
  assign _T_693 = _T_692 != 2'h0; // @[LZD.scala 39:14]
  assign _T_694 = _T_692[1]; // @[LZD.scala 39:21]
  assign _T_695 = _T_692[0]; // @[LZD.scala 39:30]
  assign _T_696 = ~ _T_695; // @[LZD.scala 39:27]
  assign _T_697 = _T_694 | _T_696; // @[LZD.scala 39:25]
  assign _T_698 = {_T_693,_T_697}; // @[Cat.scala 29:58]
  assign _T_699 = _T_691[1:0]; // @[LZD.scala 44:32]
  assign _T_700 = _T_699 != 2'h0; // @[LZD.scala 39:14]
  assign _T_701 = _T_699[1]; // @[LZD.scala 39:21]
  assign _T_702 = _T_699[0]; // @[LZD.scala 39:30]
  assign _T_703 = ~ _T_702; // @[LZD.scala 39:27]
  assign _T_704 = _T_701 | _T_703; // @[LZD.scala 39:25]
  assign _T_705 = {_T_700,_T_704}; // @[Cat.scala 29:58]
  assign _T_706 = _T_698[1]; // @[Shift.scala 12:21]
  assign _T_707 = _T_705[1]; // @[Shift.scala 12:21]
  assign _T_708 = _T_706 | _T_707; // @[LZD.scala 49:16]
  assign _T_709 = ~ _T_707; // @[LZD.scala 49:27]
  assign _T_710 = _T_706 | _T_709; // @[LZD.scala 49:25]
  assign _T_711 = _T_698[0:0]; // @[LZD.scala 49:47]
  assign _T_712 = _T_705[0:0]; // @[LZD.scala 49:59]
  assign _T_713 = _T_706 ? _T_711 : _T_712; // @[LZD.scala 49:35]
  assign _T_715 = {_T_708,_T_710,_T_713}; // @[Cat.scala 29:58]
  assign _T_716 = _T_690[3:0]; // @[LZD.scala 44:32]
  assign _T_717 = _T_716[3:2]; // @[LZD.scala 43:32]
  assign _T_718 = _T_717 != 2'h0; // @[LZD.scala 39:14]
  assign _T_719 = _T_717[1]; // @[LZD.scala 39:21]
  assign _T_720 = _T_717[0]; // @[LZD.scala 39:30]
  assign _T_721 = ~ _T_720; // @[LZD.scala 39:27]
  assign _T_722 = _T_719 | _T_721; // @[LZD.scala 39:25]
  assign _T_723 = {_T_718,_T_722}; // @[Cat.scala 29:58]
  assign _T_724 = _T_716[1:0]; // @[LZD.scala 44:32]
  assign _T_725 = _T_724 != 2'h0; // @[LZD.scala 39:14]
  assign _T_726 = _T_724[1]; // @[LZD.scala 39:21]
  assign _T_727 = _T_724[0]; // @[LZD.scala 39:30]
  assign _T_728 = ~ _T_727; // @[LZD.scala 39:27]
  assign _T_729 = _T_726 | _T_728; // @[LZD.scala 39:25]
  assign _T_730 = {_T_725,_T_729}; // @[Cat.scala 29:58]
  assign _T_731 = _T_723[1]; // @[Shift.scala 12:21]
  assign _T_732 = _T_730[1]; // @[Shift.scala 12:21]
  assign _T_733 = _T_731 | _T_732; // @[LZD.scala 49:16]
  assign _T_734 = ~ _T_732; // @[LZD.scala 49:27]
  assign _T_735 = _T_731 | _T_734; // @[LZD.scala 49:25]
  assign _T_736 = _T_723[0:0]; // @[LZD.scala 49:47]
  assign _T_737 = _T_730[0:0]; // @[LZD.scala 49:59]
  assign _T_738 = _T_731 ? _T_736 : _T_737; // @[LZD.scala 49:35]
  assign _T_740 = {_T_733,_T_735,_T_738}; // @[Cat.scala 29:58]
  assign _T_741 = _T_715[2]; // @[Shift.scala 12:21]
  assign _T_742 = _T_740[2]; // @[Shift.scala 12:21]
  assign _T_743 = _T_741 | _T_742; // @[LZD.scala 49:16]
  assign _T_744 = ~ _T_742; // @[LZD.scala 49:27]
  assign _T_745 = _T_741 | _T_744; // @[LZD.scala 49:25]
  assign _T_746 = _T_715[1:0]; // @[LZD.scala 49:47]
  assign _T_747 = _T_740[1:0]; // @[LZD.scala 49:59]
  assign _T_748 = _T_741 ? _T_746 : _T_747; // @[LZD.scala 49:35]
  assign _T_750 = {_T_743,_T_745,_T_748}; // @[Cat.scala 29:58]
  assign _T_751 = _T_689[3]; // @[Shift.scala 12:21]
  assign _T_752 = _T_750[3]; // @[Shift.scala 12:21]
  assign _T_753 = _T_751 | _T_752; // @[LZD.scala 49:16]
  assign _T_754 = ~ _T_752; // @[LZD.scala 49:27]
  assign _T_755 = _T_751 | _T_754; // @[LZD.scala 49:25]
  assign _T_756 = _T_689[2:0]; // @[LZD.scala 49:47]
  assign _T_757 = _T_750[2:0]; // @[LZD.scala 49:59]
  assign _T_758 = _T_751 ? _T_756 : _T_757; // @[LZD.scala 49:35]
  assign _T_760 = {_T_753,_T_755,_T_758}; // @[Cat.scala 29:58]
  assign _T_761 = sumXor[10:0]; // @[LZD.scala 44:32]
  assign _T_762 = _T_761[10:3]; // @[LZD.scala 43:32]
  assign _T_763 = _T_762[7:4]; // @[LZD.scala 43:32]
  assign _T_764 = _T_763[3:2]; // @[LZD.scala 43:32]
  assign _T_765 = _T_764 != 2'h0; // @[LZD.scala 39:14]
  assign _T_766 = _T_764[1]; // @[LZD.scala 39:21]
  assign _T_767 = _T_764[0]; // @[LZD.scala 39:30]
  assign _T_768 = ~ _T_767; // @[LZD.scala 39:27]
  assign _T_769 = _T_766 | _T_768; // @[LZD.scala 39:25]
  assign _T_770 = {_T_765,_T_769}; // @[Cat.scala 29:58]
  assign _T_771 = _T_763[1:0]; // @[LZD.scala 44:32]
  assign _T_772 = _T_771 != 2'h0; // @[LZD.scala 39:14]
  assign _T_773 = _T_771[1]; // @[LZD.scala 39:21]
  assign _T_774 = _T_771[0]; // @[LZD.scala 39:30]
  assign _T_775 = ~ _T_774; // @[LZD.scala 39:27]
  assign _T_776 = _T_773 | _T_775; // @[LZD.scala 39:25]
  assign _T_777 = {_T_772,_T_776}; // @[Cat.scala 29:58]
  assign _T_778 = _T_770[1]; // @[Shift.scala 12:21]
  assign _T_779 = _T_777[1]; // @[Shift.scala 12:21]
  assign _T_780 = _T_778 | _T_779; // @[LZD.scala 49:16]
  assign _T_781 = ~ _T_779; // @[LZD.scala 49:27]
  assign _T_782 = _T_778 | _T_781; // @[LZD.scala 49:25]
  assign _T_783 = _T_770[0:0]; // @[LZD.scala 49:47]
  assign _T_784 = _T_777[0:0]; // @[LZD.scala 49:59]
  assign _T_785 = _T_778 ? _T_783 : _T_784; // @[LZD.scala 49:35]
  assign _T_787 = {_T_780,_T_782,_T_785}; // @[Cat.scala 29:58]
  assign _T_788 = _T_762[3:0]; // @[LZD.scala 44:32]
  assign _T_789 = _T_788[3:2]; // @[LZD.scala 43:32]
  assign _T_790 = _T_789 != 2'h0; // @[LZD.scala 39:14]
  assign _T_791 = _T_789[1]; // @[LZD.scala 39:21]
  assign _T_792 = _T_789[0]; // @[LZD.scala 39:30]
  assign _T_793 = ~ _T_792; // @[LZD.scala 39:27]
  assign _T_794 = _T_791 | _T_793; // @[LZD.scala 39:25]
  assign _T_795 = {_T_790,_T_794}; // @[Cat.scala 29:58]
  assign _T_796 = _T_788[1:0]; // @[LZD.scala 44:32]
  assign _T_797 = _T_796 != 2'h0; // @[LZD.scala 39:14]
  assign _T_798 = _T_796[1]; // @[LZD.scala 39:21]
  assign _T_799 = _T_796[0]; // @[LZD.scala 39:30]
  assign _T_800 = ~ _T_799; // @[LZD.scala 39:27]
  assign _T_801 = _T_798 | _T_800; // @[LZD.scala 39:25]
  assign _T_802 = {_T_797,_T_801}; // @[Cat.scala 29:58]
  assign _T_803 = _T_795[1]; // @[Shift.scala 12:21]
  assign _T_804 = _T_802[1]; // @[Shift.scala 12:21]
  assign _T_805 = _T_803 | _T_804; // @[LZD.scala 49:16]
  assign _T_806 = ~ _T_804; // @[LZD.scala 49:27]
  assign _T_807 = _T_803 | _T_806; // @[LZD.scala 49:25]
  assign _T_808 = _T_795[0:0]; // @[LZD.scala 49:47]
  assign _T_809 = _T_802[0:0]; // @[LZD.scala 49:59]
  assign _T_810 = _T_803 ? _T_808 : _T_809; // @[LZD.scala 49:35]
  assign _T_812 = {_T_805,_T_807,_T_810}; // @[Cat.scala 29:58]
  assign _T_813 = _T_787[2]; // @[Shift.scala 12:21]
  assign _T_814 = _T_812[2]; // @[Shift.scala 12:21]
  assign _T_815 = _T_813 | _T_814; // @[LZD.scala 49:16]
  assign _T_816 = ~ _T_814; // @[LZD.scala 49:27]
  assign _T_817 = _T_813 | _T_816; // @[LZD.scala 49:25]
  assign _T_818 = _T_787[1:0]; // @[LZD.scala 49:47]
  assign _T_819 = _T_812[1:0]; // @[LZD.scala 49:59]
  assign _T_820 = _T_813 ? _T_818 : _T_819; // @[LZD.scala 49:35]
  assign _T_822 = {_T_815,_T_817,_T_820}; // @[Cat.scala 29:58]
  assign _T_823 = _T_761[2:0]; // @[LZD.scala 44:32]
  assign _T_824 = _T_823[2:1]; // @[LZD.scala 43:32]
  assign _T_825 = _T_824 != 2'h0; // @[LZD.scala 39:14]
  assign _T_826 = _T_824[1]; // @[LZD.scala 39:21]
  assign _T_827 = _T_824[0]; // @[LZD.scala 39:30]
  assign _T_828 = ~ _T_827; // @[LZD.scala 39:27]
  assign _T_829 = _T_826 | _T_828; // @[LZD.scala 39:25]
  assign _T_830 = {_T_825,_T_829}; // @[Cat.scala 29:58]
  assign _T_831 = _T_823[0:0]; // @[LZD.scala 44:32]
  assign _T_833 = _T_830[1]; // @[Shift.scala 12:21]
  assign _T_835 = _T_830[0:0]; // @[LZD.scala 55:32]
  assign _T_836 = _T_833 ? _T_835 : _T_831; // @[LZD.scala 55:20]
  assign _T_838 = _T_822[3]; // @[Shift.scala 12:21]
  assign _T_840 = {1'h1,_T_833,_T_836}; // @[Cat.scala 29:58]
  assign _T_841 = _T_822[2:0]; // @[LZD.scala 55:32]
  assign _T_842 = _T_838 ? _T_841 : _T_840; // @[LZD.scala 55:20]
  assign _T_843 = {_T_838,_T_842}; // @[Cat.scala 29:58]
  assign _T_844 = _T_760[4]; // @[Shift.scala 12:21]
  assign _T_846 = _T_760[3:0]; // @[LZD.scala 55:32]
  assign _T_847 = _T_844 ? _T_846 : _T_843; // @[LZD.scala 55:20]
  assign sumLZD = {_T_844,_T_847}; // @[Cat.scala 29:58]
  assign _T_848 = {1'h1,_T_844,_T_847}; // @[Cat.scala 29:58]
  assign _T_849 = $signed(_T_848); // @[PositAdder.scala 41:38]
  assign _T_851 = $signed(_T_849) + $signed(6'sh2); // @[PositAdder.scala 41:45]
  assign scaleBias = $signed(_T_851); // @[PositAdder.scala 41:45]
  assign _GEN_5 = {{3{scaleBias[5]}},scaleBias}; // @[PositAdder.scala 42:32]
  assign sumScale = $signed(greaterExp) + $signed(_GEN_5); // @[PositAdder.scala 42:32]
  assign overflow = $signed(sumScale) > $signed(10'shd0); // @[PositAdder.scala 43:30]
  assign normalShift = ~ sumLZD; // @[PositAdder.scala 44:22]
  assign _T_852 = signSumSig[25:0]; // @[PositAdder.scala 45:36]
  assign _T_853 = normalShift < 5'h1a; // @[Shift.scala 16:24]
  assign _T_855 = normalShift[4]; // @[Shift.scala 12:21]
  assign _T_856 = _T_852[9:0]; // @[Shift.scala 64:52]
  assign _T_858 = {_T_856,16'h0}; // @[Cat.scala 29:58]
  assign _T_859 = _T_855 ? _T_858 : _T_852; // @[Shift.scala 64:27]
  assign _T_860 = normalShift[3:0]; // @[Shift.scala 66:70]
  assign _T_861 = _T_860[3]; // @[Shift.scala 12:21]
  assign _T_862 = _T_859[17:0]; // @[Shift.scala 64:52]
  assign _T_864 = {_T_862,8'h0}; // @[Cat.scala 29:58]
  assign _T_865 = _T_861 ? _T_864 : _T_859; // @[Shift.scala 64:27]
  assign _T_866 = _T_860[2:0]; // @[Shift.scala 66:70]
  assign _T_867 = _T_866[2]; // @[Shift.scala 12:21]
  assign _T_868 = _T_865[21:0]; // @[Shift.scala 64:52]
  assign _T_870 = {_T_868,4'h0}; // @[Cat.scala 29:58]
  assign _T_871 = _T_867 ? _T_870 : _T_865; // @[Shift.scala 64:27]
  assign _T_872 = _T_866[1:0]; // @[Shift.scala 66:70]
  assign _T_873 = _T_872[1]; // @[Shift.scala 12:21]
  assign _T_874 = _T_871[23:0]; // @[Shift.scala 64:52]
  assign _T_876 = {_T_874,2'h0}; // @[Cat.scala 29:58]
  assign _T_877 = _T_873 ? _T_876 : _T_871; // @[Shift.scala 64:27]
  assign _T_878 = _T_872[0:0]; // @[Shift.scala 66:70]
  assign _T_880 = _T_877[24:0]; // @[Shift.scala 64:52]
  assign _T_881 = {_T_880,1'h0}; // @[Cat.scala 29:58]
  assign _T_882 = _T_878 ? _T_881 : _T_877; // @[Shift.scala 64:27]
  assign shiftSig = _T_853 ? _T_882 : 26'h0; // @[Shift.scala 16:10]
  assign _T_883 = overflow ? $signed(10'shd0) : $signed(sumScale); // @[PositAdder.scala 50:24]
  assign decS_fraction = shiftSig[25:4]; // @[PositAdder.scala 51:34]
  assign decS_isNaR = decA_isNaR | decB_isNaR; // @[PositAdder.scala 52:32]
  assign _T_886 = signSumSig != 28'h0; // @[PositAdder.scala 53:33]
  assign _T_887 = ~ _T_886; // @[PositAdder.scala 53:21]
  assign _T_888 = decA_isZero & decB_isZero; // @[PositAdder.scala 53:52]
  assign decS_isZero = _T_887 | _T_888; // @[PositAdder.scala 53:37]
  assign _T_890 = shiftSig[3:2]; // @[PositAdder.scala 54:33]
  assign _T_891 = shiftSig[1]; // @[PositAdder.scala 54:49]
  assign _T_892 = shiftSig[0]; // @[PositAdder.scala 54:63]
  assign _T_893 = _T_891 | _T_892; // @[PositAdder.scala 54:53]
  assign _GEN_6 = _T_883[8:0]; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  assign decS_scale = $signed(_GEN_6); // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  assign _T_896 = decS_scale[2:0]; // @[convert.scala 46:61]
  assign _T_897 = ~ _T_896; // @[convert.scala 46:52]
  assign _T_899 = sumSign ? _T_897 : _T_896; // @[convert.scala 46:42]
  assign _T_900 = decS_scale[8:3]; // @[convert.scala 48:34]
  assign _T_901 = _T_900[5:5]; // @[convert.scala 49:36]
  assign _T_903 = ~ _T_900; // @[convert.scala 50:36]
  assign _T_904 = $signed(_T_903); // @[convert.scala 50:36]
  assign _T_905 = _T_901 ? $signed(_T_904) : $signed(_T_900); // @[convert.scala 50:28]
  assign _T_906 = _T_901 ^ sumSign; // @[convert.scala 51:31]
  assign _T_907 = ~ _T_906; // @[convert.scala 52:43]
  assign _T_911 = {_T_907,_T_906,_T_899,decS_fraction,_T_890,_T_893}; // @[Cat.scala 29:58]
  assign _T_912 = $unsigned(_T_905); // @[Shift.scala 39:17]
  assign _T_913 = _T_912 < 6'h1e; // @[Shift.scala 39:24]
  assign _T_914 = _T_905[4:0]; // @[Shift.scala 40:44]
  assign _T_915 = _T_911[29:16]; // @[Shift.scala 90:30]
  assign _T_916 = _T_911[15:0]; // @[Shift.scala 90:48]
  assign _T_917 = _T_916 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{13'd0}, _T_917}; // @[Shift.scala 90:39]
  assign _T_918 = _T_915 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_919 = _T_914[4]; // @[Shift.scala 12:21]
  assign _T_920 = _T_911[29]; // @[Shift.scala 12:21]
  assign _T_922 = _T_920 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_923 = {_T_922,_T_918}; // @[Cat.scala 29:58]
  assign _T_924 = _T_919 ? _T_923 : _T_911; // @[Shift.scala 91:22]
  assign _T_925 = _T_914[3:0]; // @[Shift.scala 92:77]
  assign _T_926 = _T_924[29:8]; // @[Shift.scala 90:30]
  assign _T_927 = _T_924[7:0]; // @[Shift.scala 90:48]
  assign _T_928 = _T_927 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_8 = {{21'd0}, _T_928}; // @[Shift.scala 90:39]
  assign _T_929 = _T_926 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_930 = _T_925[3]; // @[Shift.scala 12:21]
  assign _T_931 = _T_924[29]; // @[Shift.scala 12:21]
  assign _T_933 = _T_931 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_934 = {_T_933,_T_929}; // @[Cat.scala 29:58]
  assign _T_935 = _T_930 ? _T_934 : _T_924; // @[Shift.scala 91:22]
  assign _T_936 = _T_925[2:0]; // @[Shift.scala 92:77]
  assign _T_937 = _T_935[29:4]; // @[Shift.scala 90:30]
  assign _T_938 = _T_935[3:0]; // @[Shift.scala 90:48]
  assign _T_939 = _T_938 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_9 = {{25'd0}, _T_939}; // @[Shift.scala 90:39]
  assign _T_940 = _T_937 | _GEN_9; // @[Shift.scala 90:39]
  assign _T_941 = _T_936[2]; // @[Shift.scala 12:21]
  assign _T_942 = _T_935[29]; // @[Shift.scala 12:21]
  assign _T_944 = _T_942 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_945 = {_T_944,_T_940}; // @[Cat.scala 29:58]
  assign _T_946 = _T_941 ? _T_945 : _T_935; // @[Shift.scala 91:22]
  assign _T_947 = _T_936[1:0]; // @[Shift.scala 92:77]
  assign _T_948 = _T_946[29:2]; // @[Shift.scala 90:30]
  assign _T_949 = _T_946[1:0]; // @[Shift.scala 90:48]
  assign _T_950 = _T_949 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_10 = {{27'd0}, _T_950}; // @[Shift.scala 90:39]
  assign _T_951 = _T_948 | _GEN_10; // @[Shift.scala 90:39]
  assign _T_952 = _T_947[1]; // @[Shift.scala 12:21]
  assign _T_953 = _T_946[29]; // @[Shift.scala 12:21]
  assign _T_955 = _T_953 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_956 = {_T_955,_T_951}; // @[Cat.scala 29:58]
  assign _T_957 = _T_952 ? _T_956 : _T_946; // @[Shift.scala 91:22]
  assign _T_958 = _T_947[0:0]; // @[Shift.scala 92:77]
  assign _T_959 = _T_957[29:1]; // @[Shift.scala 90:30]
  assign _T_960 = _T_957[0:0]; // @[Shift.scala 90:48]
  assign _GEN_11 = {{28'd0}, _T_960}; // @[Shift.scala 90:39]
  assign _T_962 = _T_959 | _GEN_11; // @[Shift.scala 90:39]
  assign _T_964 = _T_957[29]; // @[Shift.scala 12:21]
  assign _T_965 = {_T_964,_T_962}; // @[Cat.scala 29:58]
  assign _T_966 = _T_958 ? _T_965 : _T_957; // @[Shift.scala 91:22]
  assign _T_969 = _T_920 ? 30'h3fffffff : 30'h0; // @[Bitwise.scala 71:12]
  assign _T_970 = _T_913 ? _T_966 : _T_969; // @[Shift.scala 39:10]
  assign _T_971 = _T_970[3]; // @[convert.scala 55:31]
  assign _T_972 = _T_970[2]; // @[convert.scala 56:31]
  assign _T_973 = _T_970[1]; // @[convert.scala 57:31]
  assign _T_974 = _T_970[0]; // @[convert.scala 58:31]
  assign _T_975 = _T_970[29:3]; // @[convert.scala 59:69]
  assign _T_976 = _T_975 != 27'h0; // @[convert.scala 59:81]
  assign _T_977 = ~ _T_976; // @[convert.scala 59:50]
  assign _T_979 = _T_975 == 27'h7ffffff; // @[convert.scala 60:81]
  assign _T_980 = _T_971 | _T_973; // @[convert.scala 61:44]
  assign _T_981 = _T_980 | _T_974; // @[convert.scala 61:52]
  assign _T_982 = _T_972 & _T_981; // @[convert.scala 61:36]
  assign _T_983 = ~ _T_979; // @[convert.scala 62:63]
  assign _T_984 = _T_983 & _T_982; // @[convert.scala 62:103]
  assign _T_985 = _T_977 | _T_984; // @[convert.scala 62:60]
  assign _GEN_12 = {{26'd0}, _T_985}; // @[convert.scala 63:56]
  assign _T_988 = _T_975 + _GEN_12; // @[convert.scala 63:56]
  assign _T_989 = {sumSign,_T_988}; // @[Cat.scala 29:58]
  assign _T_991 = decS_isZero ? 28'h0 : _T_989; // @[Mux.scala 87:16]
  assign io_S = decS_isNaR ? 28'h8000000 : _T_991; // @[PositAdder.scala 56:8]
endmodule
