module PositMultiplier12_1(
  input         clock,
  input         reset,
  input  [11:0] io_A,
  input  [11:0] io_B,
  output [11:0] io_M
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [9:0] _T_4; // @[convert.scala 19:24]
  wire [9:0] _T_5; // @[convert.scala 19:43]
  wire [9:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [1:0] _T_68; // @[LZD.scala 44:32]
  wire  _T_69; // @[LZD.scala 39:14]
  wire  _T_70; // @[LZD.scala 39:21]
  wire  _T_71; // @[LZD.scala 39:30]
  wire  _T_72; // @[LZD.scala 39:27]
  wire  _T_73; // @[LZD.scala 39:25]
  wire  _T_75; // @[Shift.scala 12:21]
  wire [2:0] _T_77; // @[Cat.scala 29:58]
  wire [2:0] _T_78; // @[LZD.scala 55:32]
  wire [2:0] _T_79; // @[LZD.scala 55:20]
  wire [3:0] _T_80; // @[Cat.scala 29:58]
  wire [3:0] _T_81; // @[convert.scala 21:22]
  wire [8:0] _T_82; // @[convert.scala 22:36]
  wire  _T_83; // @[Shift.scala 16:24]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[Shift.scala 64:52]
  wire [8:0] _T_88; // @[Cat.scala 29:58]
  wire [8:0] _T_89; // @[Shift.scala 64:27]
  wire [2:0] _T_90; // @[Shift.scala 66:70]
  wire  _T_91; // @[Shift.scala 12:21]
  wire [4:0] _T_92; // @[Shift.scala 64:52]
  wire [8:0] _T_94; // @[Cat.scala 29:58]
  wire [8:0] _T_95; // @[Shift.scala 64:27]
  wire [1:0] _T_96; // @[Shift.scala 66:70]
  wire  _T_97; // @[Shift.scala 12:21]
  wire [6:0] _T_98; // @[Shift.scala 64:52]
  wire [8:0] _T_100; // @[Cat.scala 29:58]
  wire [8:0] _T_101; // @[Shift.scala 64:27]
  wire  _T_102; // @[Shift.scala 66:70]
  wire [7:0] _T_104; // @[Shift.scala 64:52]
  wire [8:0] _T_105; // @[Cat.scala 29:58]
  wire [8:0] _T_106; // @[Shift.scala 64:27]
  wire [8:0] _T_107; // @[Shift.scala 16:10]
  wire  _T_108; // @[convert.scala 23:34]
  wire [7:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_110; // @[convert.scala 25:26]
  wire [3:0] _T_112; // @[convert.scala 25:42]
  wire  _T_115; // @[convert.scala 26:67]
  wire  _T_116; // @[convert.scala 26:51]
  wire [5:0] _T_117; // @[Cat.scala 29:58]
  wire [10:0] _T_119; // @[convert.scala 29:56]
  wire  _T_120; // @[convert.scala 29:60]
  wire  _T_121; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_124; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_133; // @[convert.scala 18:24]
  wire  _T_134; // @[convert.scala 18:40]
  wire  _T_135; // @[convert.scala 18:36]
  wire [9:0] _T_136; // @[convert.scala 19:24]
  wire [9:0] _T_137; // @[convert.scala 19:43]
  wire [9:0] _T_138; // @[convert.scala 19:39]
  wire [7:0] _T_139; // @[LZD.scala 43:32]
  wire [3:0] _T_140; // @[LZD.scala 43:32]
  wire [1:0] _T_141; // @[LZD.scala 43:32]
  wire  _T_142; // @[LZD.scala 39:14]
  wire  _T_143; // @[LZD.scala 39:21]
  wire  _T_144; // @[LZD.scala 39:30]
  wire  _T_145; // @[LZD.scala 39:27]
  wire  _T_146; // @[LZD.scala 39:25]
  wire [1:0] _T_147; // @[Cat.scala 29:58]
  wire [1:0] _T_148; // @[LZD.scala 44:32]
  wire  _T_149; // @[LZD.scala 39:14]
  wire  _T_150; // @[LZD.scala 39:21]
  wire  _T_151; // @[LZD.scala 39:30]
  wire  _T_152; // @[LZD.scala 39:27]
  wire  _T_153; // @[LZD.scala 39:25]
  wire [1:0] _T_154; // @[Cat.scala 29:58]
  wire  _T_155; // @[Shift.scala 12:21]
  wire  _T_156; // @[Shift.scala 12:21]
  wire  _T_157; // @[LZD.scala 49:16]
  wire  _T_158; // @[LZD.scala 49:27]
  wire  _T_159; // @[LZD.scala 49:25]
  wire  _T_160; // @[LZD.scala 49:47]
  wire  _T_161; // @[LZD.scala 49:59]
  wire  _T_162; // @[LZD.scala 49:35]
  wire [2:0] _T_164; // @[Cat.scala 29:58]
  wire [3:0] _T_165; // @[LZD.scala 44:32]
  wire [1:0] _T_166; // @[LZD.scala 43:32]
  wire  _T_167; // @[LZD.scala 39:14]
  wire  _T_168; // @[LZD.scala 39:21]
  wire  _T_169; // @[LZD.scala 39:30]
  wire  _T_170; // @[LZD.scala 39:27]
  wire  _T_171; // @[LZD.scala 39:25]
  wire [1:0] _T_172; // @[Cat.scala 29:58]
  wire [1:0] _T_173; // @[LZD.scala 44:32]
  wire  _T_174; // @[LZD.scala 39:14]
  wire  _T_175; // @[LZD.scala 39:21]
  wire  _T_176; // @[LZD.scala 39:30]
  wire  _T_177; // @[LZD.scala 39:27]
  wire  _T_178; // @[LZD.scala 39:25]
  wire [1:0] _T_179; // @[Cat.scala 29:58]
  wire  _T_180; // @[Shift.scala 12:21]
  wire  _T_181; // @[Shift.scala 12:21]
  wire  _T_182; // @[LZD.scala 49:16]
  wire  _T_183; // @[LZD.scala 49:27]
  wire  _T_184; // @[LZD.scala 49:25]
  wire  _T_185; // @[LZD.scala 49:47]
  wire  _T_186; // @[LZD.scala 49:59]
  wire  _T_187; // @[LZD.scala 49:35]
  wire [2:0] _T_189; // @[Cat.scala 29:58]
  wire  _T_190; // @[Shift.scala 12:21]
  wire  _T_191; // @[Shift.scala 12:21]
  wire  _T_192; // @[LZD.scala 49:16]
  wire  _T_193; // @[LZD.scala 49:27]
  wire  _T_194; // @[LZD.scala 49:25]
  wire [1:0] _T_195; // @[LZD.scala 49:47]
  wire [1:0] _T_196; // @[LZD.scala 49:59]
  wire [1:0] _T_197; // @[LZD.scala 49:35]
  wire [3:0] _T_199; // @[Cat.scala 29:58]
  wire [1:0] _T_200; // @[LZD.scala 44:32]
  wire  _T_201; // @[LZD.scala 39:14]
  wire  _T_202; // @[LZD.scala 39:21]
  wire  _T_203; // @[LZD.scala 39:30]
  wire  _T_204; // @[LZD.scala 39:27]
  wire  _T_205; // @[LZD.scala 39:25]
  wire  _T_207; // @[Shift.scala 12:21]
  wire [2:0] _T_209; // @[Cat.scala 29:58]
  wire [2:0] _T_210; // @[LZD.scala 55:32]
  wire [2:0] _T_211; // @[LZD.scala 55:20]
  wire [3:0] _T_212; // @[Cat.scala 29:58]
  wire [3:0] _T_213; // @[convert.scala 21:22]
  wire [8:0] _T_214; // @[convert.scala 22:36]
  wire  _T_215; // @[Shift.scala 16:24]
  wire  _T_217; // @[Shift.scala 12:21]
  wire  _T_218; // @[Shift.scala 64:52]
  wire [8:0] _T_220; // @[Cat.scala 29:58]
  wire [8:0] _T_221; // @[Shift.scala 64:27]
  wire [2:0] _T_222; // @[Shift.scala 66:70]
  wire  _T_223; // @[Shift.scala 12:21]
  wire [4:0] _T_224; // @[Shift.scala 64:52]
  wire [8:0] _T_226; // @[Cat.scala 29:58]
  wire [8:0] _T_227; // @[Shift.scala 64:27]
  wire [1:0] _T_228; // @[Shift.scala 66:70]
  wire  _T_229; // @[Shift.scala 12:21]
  wire [6:0] _T_230; // @[Shift.scala 64:52]
  wire [8:0] _T_232; // @[Cat.scala 29:58]
  wire [8:0] _T_233; // @[Shift.scala 64:27]
  wire  _T_234; // @[Shift.scala 66:70]
  wire [7:0] _T_236; // @[Shift.scala 64:52]
  wire [8:0] _T_237; // @[Cat.scala 29:58]
  wire [8:0] _T_238; // @[Shift.scala 64:27]
  wire [8:0] _T_239; // @[Shift.scala 16:10]
  wire  _T_240; // @[convert.scala 23:34]
  wire [7:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_242; // @[convert.scala 25:26]
  wire [3:0] _T_244; // @[convert.scala 25:42]
  wire  _T_247; // @[convert.scala 26:67]
  wire  _T_248; // @[convert.scala 26:51]
  wire [5:0] _T_249; // @[Cat.scala 29:58]
  wire [10:0] _T_251; // @[convert.scala 29:56]
  wire  _T_252; // @[convert.scala 29:60]
  wire  _T_253; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_256; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_264; // @[PositMultiplier.scala 43:34]
  wire [9:0] _T_266; // @[Cat.scala 29:58]
  wire [9:0] sigA; // @[PositMultiplier.scala 43:61]
  wire  _T_267; // @[PositMultiplier.scala 44:34]
  wire [9:0] _T_269; // @[Cat.scala 29:58]
  wire [9:0] sigB; // @[PositMultiplier.scala 44:61]
  wire [19:0] _T_270; // @[PositMultiplier.scala 45:25]
  wire [19:0] sigP; // @[PositMultiplier.scala 45:33]
  wire [1:0] head2; // @[PositMultiplier.scala 46:28]
  wire  _T_271; // @[PositMultiplier.scala 47:31]
  wire  _T_272; // @[PositMultiplier.scala 47:25]
  wire  _T_273; // @[PositMultiplier.scala 47:42]
  wire  addTwo; // @[PositMultiplier.scala 47:35]
  wire  _T_274; // @[PositMultiplier.scala 49:23]
  wire  _T_275; // @[PositMultiplier.scala 49:49]
  wire  addOne; // @[PositMultiplier.scala 49:43]
  wire [1:0] _T_276; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositMultiplier.scala 50:39]
  wire [16:0] _T_277; // @[PositMultiplier.scala 53:81]
  wire [15:0] _T_278; // @[PositMultiplier.scala 54:81]
  wire [16:0] _T_279; // @[PositMultiplier.scala 54:104]
  wire [16:0] frac; // @[PositMultiplier.scala 51:22]
  wire [6:0] _T_280; // @[PositMultiplier.scala 56:30]
  wire [6:0] _GEN_0; // @[PositMultiplier.scala 56:44]
  wire [6:0] _T_282; // @[PositMultiplier.scala 56:44]
  wire [6:0] mulScale; // @[PositMultiplier.scala 56:44]
  wire  underflow; // @[PositMultiplier.scala 57:28]
  wire  overflow; // @[PositMultiplier.scala 58:28]
  wire  decM_sign; // @[PositMultiplier.scala 62:29]
  wire [6:0] _T_285; // @[Mux.scala 87:16]
  wire [6:0] _T_286; // @[Mux.scala 87:16]
  wire [7:0] decM_fraction; // @[PositMultiplier.scala 70:29]
  wire  decM_isNaR; // @[PositMultiplier.scala 71:31]
  wire  decM_isZero; // @[PositMultiplier.scala 72:32]
  wire [8:0] grsTmp; // @[PositMultiplier.scala 75:30]
  wire [1:0] _T_290; // @[PositMultiplier.scala 78:32]
  wire [6:0] _T_291; // @[PositMultiplier.scala 78:48]
  wire  _T_292; // @[PositMultiplier.scala 78:52]
  wire [5:0] _GEN_1; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  wire [5:0] decM_scale; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  wire  _T_295; // @[convert.scala 46:61]
  wire  _T_296; // @[convert.scala 46:52]
  wire  _T_298; // @[convert.scala 46:42]
  wire [4:0] _T_299; // @[convert.scala 48:34]
  wire  _T_300; // @[convert.scala 49:36]
  wire [4:0] _T_302; // @[convert.scala 50:36]
  wire [4:0] _T_303; // @[convert.scala 50:36]
  wire [4:0] _T_304; // @[convert.scala 50:28]
  wire  _T_305; // @[convert.scala 51:31]
  wire  _T_306; // @[convert.scala 52:43]
  wire [13:0] _T_310; // @[Cat.scala 29:58]
  wire [4:0] _T_311; // @[Shift.scala 39:17]
  wire  _T_312; // @[Shift.scala 39:24]
  wire [3:0] _T_313; // @[Shift.scala 40:44]
  wire [5:0] _T_314; // @[Shift.scala 90:30]
  wire [7:0] _T_315; // @[Shift.scala 90:48]
  wire  _T_316; // @[Shift.scala 90:57]
  wire [5:0] _GEN_2; // @[Shift.scala 90:39]
  wire [5:0] _T_317; // @[Shift.scala 90:39]
  wire  _T_318; // @[Shift.scala 12:21]
  wire  _T_319; // @[Shift.scala 12:21]
  wire [7:0] _T_321; // @[Bitwise.scala 71:12]
  wire [13:0] _T_322; // @[Cat.scala 29:58]
  wire [13:0] _T_323; // @[Shift.scala 91:22]
  wire [2:0] _T_324; // @[Shift.scala 92:77]
  wire [9:0] _T_325; // @[Shift.scala 90:30]
  wire [3:0] _T_326; // @[Shift.scala 90:48]
  wire  _T_327; // @[Shift.scala 90:57]
  wire [9:0] _GEN_3; // @[Shift.scala 90:39]
  wire [9:0] _T_328; // @[Shift.scala 90:39]
  wire  _T_329; // @[Shift.scala 12:21]
  wire  _T_330; // @[Shift.scala 12:21]
  wire [3:0] _T_332; // @[Bitwise.scala 71:12]
  wire [13:0] _T_333; // @[Cat.scala 29:58]
  wire [13:0] _T_334; // @[Shift.scala 91:22]
  wire [1:0] _T_335; // @[Shift.scala 92:77]
  wire [11:0] _T_336; // @[Shift.scala 90:30]
  wire [1:0] _T_337; // @[Shift.scala 90:48]
  wire  _T_338; // @[Shift.scala 90:57]
  wire [11:0] _GEN_4; // @[Shift.scala 90:39]
  wire [11:0] _T_339; // @[Shift.scala 90:39]
  wire  _T_340; // @[Shift.scala 12:21]
  wire  _T_341; // @[Shift.scala 12:21]
  wire [1:0] _T_343; // @[Bitwise.scala 71:12]
  wire [13:0] _T_344; // @[Cat.scala 29:58]
  wire [13:0] _T_345; // @[Shift.scala 91:22]
  wire  _T_346; // @[Shift.scala 92:77]
  wire [12:0] _T_347; // @[Shift.scala 90:30]
  wire  _T_348; // @[Shift.scala 90:48]
  wire [12:0] _GEN_5; // @[Shift.scala 90:39]
  wire [12:0] _T_350; // @[Shift.scala 90:39]
  wire  _T_352; // @[Shift.scala 12:21]
  wire [13:0] _T_353; // @[Cat.scala 29:58]
  wire [13:0] _T_354; // @[Shift.scala 91:22]
  wire [13:0] _T_357; // @[Bitwise.scala 71:12]
  wire [13:0] _T_358; // @[Shift.scala 39:10]
  wire  _T_359; // @[convert.scala 55:31]
  wire  _T_360; // @[convert.scala 56:31]
  wire  _T_361; // @[convert.scala 57:31]
  wire  _T_362; // @[convert.scala 58:31]
  wire [10:0] _T_363; // @[convert.scala 59:69]
  wire  _T_364; // @[convert.scala 59:81]
  wire  _T_365; // @[convert.scala 59:50]
  wire  _T_367; // @[convert.scala 60:81]
  wire  _T_368; // @[convert.scala 61:44]
  wire  _T_369; // @[convert.scala 61:52]
  wire  _T_370; // @[convert.scala 61:36]
  wire  _T_371; // @[convert.scala 62:63]
  wire  _T_372; // @[convert.scala 62:103]
  wire  _T_373; // @[convert.scala 62:60]
  wire [10:0] _GEN_6; // @[convert.scala 63:56]
  wire [10:0] _T_376; // @[convert.scala 63:56]
  wire [11:0] _T_377; // @[Cat.scala 29:58]
  wire [11:0] _T_379; // @[Mux.scala 87:16]
  assign _T_1 = io_A[11]; // @[convert.scala 18:24]
  assign _T_2 = io_A[10]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[10:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[9:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[9:2]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[1:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68 != 2'h0; // @[LZD.scala 39:14]
  assign _T_70 = _T_68[1]; // @[LZD.scala 39:21]
  assign _T_71 = _T_68[0]; // @[LZD.scala 39:30]
  assign _T_72 = ~ _T_71; // @[LZD.scala 39:27]
  assign _T_73 = _T_70 | _T_72; // @[LZD.scala 39:25]
  assign _T_75 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_77 = {1'h1,_T_69,_T_73}; // @[Cat.scala 29:58]
  assign _T_78 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_79 = _T_75 ? _T_78 : _T_77; // @[LZD.scala 55:20]
  assign _T_80 = {_T_75,_T_79}; // @[Cat.scala 29:58]
  assign _T_81 = ~ _T_80; // @[convert.scala 21:22]
  assign _T_82 = io_A[8:0]; // @[convert.scala 22:36]
  assign _T_83 = _T_81 < 4'h9; // @[Shift.scala 16:24]
  assign _T_85 = _T_81[3]; // @[Shift.scala 12:21]
  assign _T_86 = _T_82[0:0]; // @[Shift.scala 64:52]
  assign _T_88 = {_T_86,8'h0}; // @[Cat.scala 29:58]
  assign _T_89 = _T_85 ? _T_88 : _T_82; // @[Shift.scala 64:27]
  assign _T_90 = _T_81[2:0]; // @[Shift.scala 66:70]
  assign _T_91 = _T_90[2]; // @[Shift.scala 12:21]
  assign _T_92 = _T_89[4:0]; // @[Shift.scala 64:52]
  assign _T_94 = {_T_92,4'h0}; // @[Cat.scala 29:58]
  assign _T_95 = _T_91 ? _T_94 : _T_89; // @[Shift.scala 64:27]
  assign _T_96 = _T_90[1:0]; // @[Shift.scala 66:70]
  assign _T_97 = _T_96[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_95[6:0]; // @[Shift.scala 64:52]
  assign _T_100 = {_T_98,2'h0}; // @[Cat.scala 29:58]
  assign _T_101 = _T_97 ? _T_100 : _T_95; // @[Shift.scala 64:27]
  assign _T_102 = _T_96[0:0]; // @[Shift.scala 66:70]
  assign _T_104 = _T_101[7:0]; // @[Shift.scala 64:52]
  assign _T_105 = {_T_104,1'h0}; // @[Cat.scala 29:58]
  assign _T_106 = _T_102 ? _T_105 : _T_101; // @[Shift.scala 64:27]
  assign _T_107 = _T_83 ? _T_106 : 9'h0; // @[Shift.scala 16:10]
  assign _T_108 = _T_107[8:8]; // @[convert.scala 23:34]
  assign decA_fraction = _T_107[7:0]; // @[convert.scala 24:34]
  assign _T_110 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_112 = _T_3 ? _T_81 : _T_80; // @[convert.scala 25:42]
  assign _T_115 = ~ _T_108; // @[convert.scala 26:67]
  assign _T_116 = _T_1 ? _T_115 : _T_108; // @[convert.scala 26:51]
  assign _T_117 = {_T_110,_T_112,_T_116}; // @[Cat.scala 29:58]
  assign _T_119 = io_A[10:0]; // @[convert.scala 29:56]
  assign _T_120 = _T_119 != 11'h0; // @[convert.scala 29:60]
  assign _T_121 = ~ _T_120; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_121; // @[convert.scala 29:39]
  assign _T_124 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_124 & _T_121; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_117); // @[convert.scala 32:24]
  assign _T_133 = io_B[11]; // @[convert.scala 18:24]
  assign _T_134 = io_B[10]; // @[convert.scala 18:40]
  assign _T_135 = _T_133 ^ _T_134; // @[convert.scala 18:36]
  assign _T_136 = io_B[10:1]; // @[convert.scala 19:24]
  assign _T_137 = io_B[9:0]; // @[convert.scala 19:43]
  assign _T_138 = _T_136 ^ _T_137; // @[convert.scala 19:39]
  assign _T_139 = _T_138[9:2]; // @[LZD.scala 43:32]
  assign _T_140 = _T_139[7:4]; // @[LZD.scala 43:32]
  assign _T_141 = _T_140[3:2]; // @[LZD.scala 43:32]
  assign _T_142 = _T_141 != 2'h0; // @[LZD.scala 39:14]
  assign _T_143 = _T_141[1]; // @[LZD.scala 39:21]
  assign _T_144 = _T_141[0]; // @[LZD.scala 39:30]
  assign _T_145 = ~ _T_144; // @[LZD.scala 39:27]
  assign _T_146 = _T_143 | _T_145; // @[LZD.scala 39:25]
  assign _T_147 = {_T_142,_T_146}; // @[Cat.scala 29:58]
  assign _T_148 = _T_140[1:0]; // @[LZD.scala 44:32]
  assign _T_149 = _T_148 != 2'h0; // @[LZD.scala 39:14]
  assign _T_150 = _T_148[1]; // @[LZD.scala 39:21]
  assign _T_151 = _T_148[0]; // @[LZD.scala 39:30]
  assign _T_152 = ~ _T_151; // @[LZD.scala 39:27]
  assign _T_153 = _T_150 | _T_152; // @[LZD.scala 39:25]
  assign _T_154 = {_T_149,_T_153}; // @[Cat.scala 29:58]
  assign _T_155 = _T_147[1]; // @[Shift.scala 12:21]
  assign _T_156 = _T_154[1]; // @[Shift.scala 12:21]
  assign _T_157 = _T_155 | _T_156; // @[LZD.scala 49:16]
  assign _T_158 = ~ _T_156; // @[LZD.scala 49:27]
  assign _T_159 = _T_155 | _T_158; // @[LZD.scala 49:25]
  assign _T_160 = _T_147[0:0]; // @[LZD.scala 49:47]
  assign _T_161 = _T_154[0:0]; // @[LZD.scala 49:59]
  assign _T_162 = _T_155 ? _T_160 : _T_161; // @[LZD.scala 49:35]
  assign _T_164 = {_T_157,_T_159,_T_162}; // @[Cat.scala 29:58]
  assign _T_165 = _T_139[3:0]; // @[LZD.scala 44:32]
  assign _T_166 = _T_165[3:2]; // @[LZD.scala 43:32]
  assign _T_167 = _T_166 != 2'h0; // @[LZD.scala 39:14]
  assign _T_168 = _T_166[1]; // @[LZD.scala 39:21]
  assign _T_169 = _T_166[0]; // @[LZD.scala 39:30]
  assign _T_170 = ~ _T_169; // @[LZD.scala 39:27]
  assign _T_171 = _T_168 | _T_170; // @[LZD.scala 39:25]
  assign _T_172 = {_T_167,_T_171}; // @[Cat.scala 29:58]
  assign _T_173 = _T_165[1:0]; // @[LZD.scala 44:32]
  assign _T_174 = _T_173 != 2'h0; // @[LZD.scala 39:14]
  assign _T_175 = _T_173[1]; // @[LZD.scala 39:21]
  assign _T_176 = _T_173[0]; // @[LZD.scala 39:30]
  assign _T_177 = ~ _T_176; // @[LZD.scala 39:27]
  assign _T_178 = _T_175 | _T_177; // @[LZD.scala 39:25]
  assign _T_179 = {_T_174,_T_178}; // @[Cat.scala 29:58]
  assign _T_180 = _T_172[1]; // @[Shift.scala 12:21]
  assign _T_181 = _T_179[1]; // @[Shift.scala 12:21]
  assign _T_182 = _T_180 | _T_181; // @[LZD.scala 49:16]
  assign _T_183 = ~ _T_181; // @[LZD.scala 49:27]
  assign _T_184 = _T_180 | _T_183; // @[LZD.scala 49:25]
  assign _T_185 = _T_172[0:0]; // @[LZD.scala 49:47]
  assign _T_186 = _T_179[0:0]; // @[LZD.scala 49:59]
  assign _T_187 = _T_180 ? _T_185 : _T_186; // @[LZD.scala 49:35]
  assign _T_189 = {_T_182,_T_184,_T_187}; // @[Cat.scala 29:58]
  assign _T_190 = _T_164[2]; // @[Shift.scala 12:21]
  assign _T_191 = _T_189[2]; // @[Shift.scala 12:21]
  assign _T_192 = _T_190 | _T_191; // @[LZD.scala 49:16]
  assign _T_193 = ~ _T_191; // @[LZD.scala 49:27]
  assign _T_194 = _T_190 | _T_193; // @[LZD.scala 49:25]
  assign _T_195 = _T_164[1:0]; // @[LZD.scala 49:47]
  assign _T_196 = _T_189[1:0]; // @[LZD.scala 49:59]
  assign _T_197 = _T_190 ? _T_195 : _T_196; // @[LZD.scala 49:35]
  assign _T_199 = {_T_192,_T_194,_T_197}; // @[Cat.scala 29:58]
  assign _T_200 = _T_138[1:0]; // @[LZD.scala 44:32]
  assign _T_201 = _T_200 != 2'h0; // @[LZD.scala 39:14]
  assign _T_202 = _T_200[1]; // @[LZD.scala 39:21]
  assign _T_203 = _T_200[0]; // @[LZD.scala 39:30]
  assign _T_204 = ~ _T_203; // @[LZD.scala 39:27]
  assign _T_205 = _T_202 | _T_204; // @[LZD.scala 39:25]
  assign _T_207 = _T_199[3]; // @[Shift.scala 12:21]
  assign _T_209 = {1'h1,_T_201,_T_205}; // @[Cat.scala 29:58]
  assign _T_210 = _T_199[2:0]; // @[LZD.scala 55:32]
  assign _T_211 = _T_207 ? _T_210 : _T_209; // @[LZD.scala 55:20]
  assign _T_212 = {_T_207,_T_211}; // @[Cat.scala 29:58]
  assign _T_213 = ~ _T_212; // @[convert.scala 21:22]
  assign _T_214 = io_B[8:0]; // @[convert.scala 22:36]
  assign _T_215 = _T_213 < 4'h9; // @[Shift.scala 16:24]
  assign _T_217 = _T_213[3]; // @[Shift.scala 12:21]
  assign _T_218 = _T_214[0:0]; // @[Shift.scala 64:52]
  assign _T_220 = {_T_218,8'h0}; // @[Cat.scala 29:58]
  assign _T_221 = _T_217 ? _T_220 : _T_214; // @[Shift.scala 64:27]
  assign _T_222 = _T_213[2:0]; // @[Shift.scala 66:70]
  assign _T_223 = _T_222[2]; // @[Shift.scala 12:21]
  assign _T_224 = _T_221[4:0]; // @[Shift.scala 64:52]
  assign _T_226 = {_T_224,4'h0}; // @[Cat.scala 29:58]
  assign _T_227 = _T_223 ? _T_226 : _T_221; // @[Shift.scala 64:27]
  assign _T_228 = _T_222[1:0]; // @[Shift.scala 66:70]
  assign _T_229 = _T_228[1]; // @[Shift.scala 12:21]
  assign _T_230 = _T_227[6:0]; // @[Shift.scala 64:52]
  assign _T_232 = {_T_230,2'h0}; // @[Cat.scala 29:58]
  assign _T_233 = _T_229 ? _T_232 : _T_227; // @[Shift.scala 64:27]
  assign _T_234 = _T_228[0:0]; // @[Shift.scala 66:70]
  assign _T_236 = _T_233[7:0]; // @[Shift.scala 64:52]
  assign _T_237 = {_T_236,1'h0}; // @[Cat.scala 29:58]
  assign _T_238 = _T_234 ? _T_237 : _T_233; // @[Shift.scala 64:27]
  assign _T_239 = _T_215 ? _T_238 : 9'h0; // @[Shift.scala 16:10]
  assign _T_240 = _T_239[8:8]; // @[convert.scala 23:34]
  assign decB_fraction = _T_239[7:0]; // @[convert.scala 24:34]
  assign _T_242 = _T_135 == 1'h0; // @[convert.scala 25:26]
  assign _T_244 = _T_135 ? _T_213 : _T_212; // @[convert.scala 25:42]
  assign _T_247 = ~ _T_240; // @[convert.scala 26:67]
  assign _T_248 = _T_133 ? _T_247 : _T_240; // @[convert.scala 26:51]
  assign _T_249 = {_T_242,_T_244,_T_248}; // @[Cat.scala 29:58]
  assign _T_251 = io_B[10:0]; // @[convert.scala 29:56]
  assign _T_252 = _T_251 != 11'h0; // @[convert.scala 29:60]
  assign _T_253 = ~ _T_252; // @[convert.scala 29:41]
  assign decB_isNaR = _T_133 & _T_253; // @[convert.scala 29:39]
  assign _T_256 = _T_133 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_256 & _T_253; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_249); // @[convert.scala 32:24]
  assign _T_264 = ~ _T_1; // @[PositMultiplier.scala 43:34]
  assign _T_266 = {_T_1,_T_264,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_266); // @[PositMultiplier.scala 43:61]
  assign _T_267 = ~ _T_133; // @[PositMultiplier.scala 44:34]
  assign _T_269 = {_T_133,_T_267,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_269); // @[PositMultiplier.scala 44:61]
  assign _T_270 = $signed(sigA) * $signed(sigB); // @[PositMultiplier.scala 45:25]
  assign sigP = $unsigned(_T_270); // @[PositMultiplier.scala 45:33]
  assign head2 = sigP[19:18]; // @[PositMultiplier.scala 46:28]
  assign _T_271 = head2[1]; // @[PositMultiplier.scala 47:31]
  assign _T_272 = ~ _T_271; // @[PositMultiplier.scala 47:25]
  assign _T_273 = head2[0]; // @[PositMultiplier.scala 47:42]
  assign addTwo = _T_272 & _T_273; // @[PositMultiplier.scala 47:35]
  assign _T_274 = sigP[19]; // @[PositMultiplier.scala 49:23]
  assign _T_275 = sigP[17]; // @[PositMultiplier.scala 49:49]
  assign addOne = _T_274 ^ _T_275; // @[PositMultiplier.scala 49:43]
  assign _T_276 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_276)}; // @[PositMultiplier.scala 50:39]
  assign _T_277 = sigP[16:0]; // @[PositMultiplier.scala 53:81]
  assign _T_278 = sigP[15:0]; // @[PositMultiplier.scala 54:81]
  assign _T_279 = {_T_278, 1'h0}; // @[PositMultiplier.scala 54:104]
  assign frac = addOne ? _T_277 : _T_279; // @[PositMultiplier.scala 51:22]
  assign _T_280 = $signed(decA_scale) + $signed(decB_scale); // @[PositMultiplier.scala 56:30]
  assign _GEN_0 = {{4{expBias[2]}},expBias}; // @[PositMultiplier.scala 56:44]
  assign _T_282 = $signed(_T_280) + $signed(_GEN_0); // @[PositMultiplier.scala 56:44]
  assign mulScale = $signed(_T_282); // @[PositMultiplier.scala 56:44]
  assign underflow = $signed(mulScale) < $signed(-7'sh14); // @[PositMultiplier.scala 57:28]
  assign overflow = $signed(mulScale) > $signed(7'sh14); // @[PositMultiplier.scala 58:28]
  assign decM_sign = sigP[19:19]; // @[PositMultiplier.scala 62:29]
  assign _T_285 = underflow ? $signed(-7'sh14) : $signed(mulScale); // @[Mux.scala 87:16]
  assign _T_286 = overflow ? $signed(7'sh14) : $signed(_T_285); // @[Mux.scala 87:16]
  assign decM_fraction = frac[16:9]; // @[PositMultiplier.scala 70:29]
  assign decM_isNaR = decA_isNaR | decB_isNaR; // @[PositMultiplier.scala 71:31]
  assign decM_isZero = decA_isZero | decB_isZero; // @[PositMultiplier.scala 72:32]
  assign grsTmp = frac[8:0]; // @[PositMultiplier.scala 75:30]
  assign _T_290 = grsTmp[8:7]; // @[PositMultiplier.scala 78:32]
  assign _T_291 = grsTmp[6:0]; // @[PositMultiplier.scala 78:48]
  assign _T_292 = _T_291 != 7'h0; // @[PositMultiplier.scala 78:52]
  assign _GEN_1 = _T_286[5:0]; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  assign decM_scale = $signed(_GEN_1); // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  assign _T_295 = decM_scale[0]; // @[convert.scala 46:61]
  assign _T_296 = ~ _T_295; // @[convert.scala 46:52]
  assign _T_298 = decM_sign ? _T_296 : _T_295; // @[convert.scala 46:42]
  assign _T_299 = decM_scale[5:1]; // @[convert.scala 48:34]
  assign _T_300 = _T_299[4:4]; // @[convert.scala 49:36]
  assign _T_302 = ~ _T_299; // @[convert.scala 50:36]
  assign _T_303 = $signed(_T_302); // @[convert.scala 50:36]
  assign _T_304 = _T_300 ? $signed(_T_303) : $signed(_T_299); // @[convert.scala 50:28]
  assign _T_305 = _T_300 ^ decM_sign; // @[convert.scala 51:31]
  assign _T_306 = ~ _T_305; // @[convert.scala 52:43]
  assign _T_310 = {_T_306,_T_305,_T_298,decM_fraction,_T_290,_T_292}; // @[Cat.scala 29:58]
  assign _T_311 = $unsigned(_T_304); // @[Shift.scala 39:17]
  assign _T_312 = _T_311 < 5'he; // @[Shift.scala 39:24]
  assign _T_313 = _T_304[3:0]; // @[Shift.scala 40:44]
  assign _T_314 = _T_310[13:8]; // @[Shift.scala 90:30]
  assign _T_315 = _T_310[7:0]; // @[Shift.scala 90:48]
  assign _T_316 = _T_315 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{5'd0}, _T_316}; // @[Shift.scala 90:39]
  assign _T_317 = _T_314 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_318 = _T_313[3]; // @[Shift.scala 12:21]
  assign _T_319 = _T_310[13]; // @[Shift.scala 12:21]
  assign _T_321 = _T_319 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_322 = {_T_321,_T_317}; // @[Cat.scala 29:58]
  assign _T_323 = _T_318 ? _T_322 : _T_310; // @[Shift.scala 91:22]
  assign _T_324 = _T_313[2:0]; // @[Shift.scala 92:77]
  assign _T_325 = _T_323[13:4]; // @[Shift.scala 90:30]
  assign _T_326 = _T_323[3:0]; // @[Shift.scala 90:48]
  assign _T_327 = _T_326 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_3 = {{9'd0}, _T_327}; // @[Shift.scala 90:39]
  assign _T_328 = _T_325 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_329 = _T_324[2]; // @[Shift.scala 12:21]
  assign _T_330 = _T_323[13]; // @[Shift.scala 12:21]
  assign _T_332 = _T_330 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_333 = {_T_332,_T_328}; // @[Cat.scala 29:58]
  assign _T_334 = _T_329 ? _T_333 : _T_323; // @[Shift.scala 91:22]
  assign _T_335 = _T_324[1:0]; // @[Shift.scala 92:77]
  assign _T_336 = _T_334[13:2]; // @[Shift.scala 90:30]
  assign _T_337 = _T_334[1:0]; // @[Shift.scala 90:48]
  assign _T_338 = _T_337 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_4 = {{11'd0}, _T_338}; // @[Shift.scala 90:39]
  assign _T_339 = _T_336 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_340 = _T_335[1]; // @[Shift.scala 12:21]
  assign _T_341 = _T_334[13]; // @[Shift.scala 12:21]
  assign _T_343 = _T_341 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_344 = {_T_343,_T_339}; // @[Cat.scala 29:58]
  assign _T_345 = _T_340 ? _T_344 : _T_334; // @[Shift.scala 91:22]
  assign _T_346 = _T_335[0:0]; // @[Shift.scala 92:77]
  assign _T_347 = _T_345[13:1]; // @[Shift.scala 90:30]
  assign _T_348 = _T_345[0:0]; // @[Shift.scala 90:48]
  assign _GEN_5 = {{12'd0}, _T_348}; // @[Shift.scala 90:39]
  assign _T_350 = _T_347 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_352 = _T_345[13]; // @[Shift.scala 12:21]
  assign _T_353 = {_T_352,_T_350}; // @[Cat.scala 29:58]
  assign _T_354 = _T_346 ? _T_353 : _T_345; // @[Shift.scala 91:22]
  assign _T_357 = _T_319 ? 14'h3fff : 14'h0; // @[Bitwise.scala 71:12]
  assign _T_358 = _T_312 ? _T_354 : _T_357; // @[Shift.scala 39:10]
  assign _T_359 = _T_358[3]; // @[convert.scala 55:31]
  assign _T_360 = _T_358[2]; // @[convert.scala 56:31]
  assign _T_361 = _T_358[1]; // @[convert.scala 57:31]
  assign _T_362 = _T_358[0]; // @[convert.scala 58:31]
  assign _T_363 = _T_358[13:3]; // @[convert.scala 59:69]
  assign _T_364 = _T_363 != 11'h0; // @[convert.scala 59:81]
  assign _T_365 = ~ _T_364; // @[convert.scala 59:50]
  assign _T_367 = _T_363 == 11'h7ff; // @[convert.scala 60:81]
  assign _T_368 = _T_359 | _T_361; // @[convert.scala 61:44]
  assign _T_369 = _T_368 | _T_362; // @[convert.scala 61:52]
  assign _T_370 = _T_360 & _T_369; // @[convert.scala 61:36]
  assign _T_371 = ~ _T_367; // @[convert.scala 62:63]
  assign _T_372 = _T_371 & _T_370; // @[convert.scala 62:103]
  assign _T_373 = _T_365 | _T_372; // @[convert.scala 62:60]
  assign _GEN_6 = {{10'd0}, _T_373}; // @[convert.scala 63:56]
  assign _T_376 = _T_363 + _GEN_6; // @[convert.scala 63:56]
  assign _T_377 = {decM_sign,_T_376}; // @[Cat.scala 29:58]
  assign _T_379 = decM_isZero ? 12'h0 : _T_377; // @[Mux.scala 87:16]
  assign io_M = decM_isNaR ? 12'h800 : _T_379; // @[PositMultiplier.scala 86:8]
endmodule
