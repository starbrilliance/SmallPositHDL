module PositFMA12_1(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [1:0]  io_fmaOp,
  input  [11:0] io_A,
  input  [11:0] io_B,
  input  [11:0] io_C,
  output [11:0] io_F,
  output        io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [11:0] _T_2; // @[Bitwise.scala 71:12]
  wire [11:0] _T_3; // @[PositFMA.scala 47:41]
  wire [11:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [11:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [11:0] _T_8; // @[Bitwise.scala 71:12]
  wire [11:0] _T_9; // @[PositFMA.scala 48:41]
  wire [11:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [11:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [9:0] _T_16; // @[convert.scala 19:24]
  wire [9:0] _T_17; // @[convert.scala 19:43]
  wire [9:0] _T_18; // @[convert.scala 19:39]
  wire [7:0] _T_19; // @[LZD.scala 43:32]
  wire [3:0] _T_20; // @[LZD.scala 43:32]
  wire [1:0] _T_21; // @[LZD.scala 43:32]
  wire  _T_22; // @[LZD.scala 39:14]
  wire  _T_23; // @[LZD.scala 39:21]
  wire  _T_24; // @[LZD.scala 39:30]
  wire  _T_25; // @[LZD.scala 39:27]
  wire  _T_26; // @[LZD.scala 39:25]
  wire [1:0] _T_27; // @[Cat.scala 29:58]
  wire [1:0] _T_28; // @[LZD.scala 44:32]
  wire  _T_29; // @[LZD.scala 39:14]
  wire  _T_30; // @[LZD.scala 39:21]
  wire  _T_31; // @[LZD.scala 39:30]
  wire  _T_32; // @[LZD.scala 39:27]
  wire  _T_33; // @[LZD.scala 39:25]
  wire [1:0] _T_34; // @[Cat.scala 29:58]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[Shift.scala 12:21]
  wire  _T_37; // @[LZD.scala 49:16]
  wire  _T_38; // @[LZD.scala 49:27]
  wire  _T_39; // @[LZD.scala 49:25]
  wire  _T_40; // @[LZD.scala 49:47]
  wire  _T_41; // @[LZD.scala 49:59]
  wire  _T_42; // @[LZD.scala 49:35]
  wire [2:0] _T_44; // @[Cat.scala 29:58]
  wire [3:0] _T_45; // @[LZD.scala 44:32]
  wire [1:0] _T_46; // @[LZD.scala 43:32]
  wire  _T_47; // @[LZD.scala 39:14]
  wire  _T_48; // @[LZD.scala 39:21]
  wire  _T_49; // @[LZD.scala 39:30]
  wire  _T_50; // @[LZD.scala 39:27]
  wire  _T_51; // @[LZD.scala 39:25]
  wire [1:0] _T_52; // @[Cat.scala 29:58]
  wire [1:0] _T_53; // @[LZD.scala 44:32]
  wire  _T_54; // @[LZD.scala 39:14]
  wire  _T_55; // @[LZD.scala 39:21]
  wire  _T_56; // @[LZD.scala 39:30]
  wire  _T_57; // @[LZD.scala 39:27]
  wire  _T_58; // @[LZD.scala 39:25]
  wire [1:0] _T_59; // @[Cat.scala 29:58]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[LZD.scala 49:16]
  wire  _T_63; // @[LZD.scala 49:27]
  wire  _T_64; // @[LZD.scala 49:25]
  wire  _T_65; // @[LZD.scala 49:47]
  wire  _T_66; // @[LZD.scala 49:59]
  wire  _T_67; // @[LZD.scala 49:35]
  wire [2:0] _T_69; // @[Cat.scala 29:58]
  wire  _T_70; // @[Shift.scala 12:21]
  wire  _T_71; // @[Shift.scala 12:21]
  wire  _T_72; // @[LZD.scala 49:16]
  wire  _T_73; // @[LZD.scala 49:27]
  wire  _T_74; // @[LZD.scala 49:25]
  wire [1:0] _T_75; // @[LZD.scala 49:47]
  wire [1:0] _T_76; // @[LZD.scala 49:59]
  wire [1:0] _T_77; // @[LZD.scala 49:35]
  wire [3:0] _T_79; // @[Cat.scala 29:58]
  wire [1:0] _T_80; // @[LZD.scala 44:32]
  wire  _T_81; // @[LZD.scala 39:14]
  wire  _T_82; // @[LZD.scala 39:21]
  wire  _T_83; // @[LZD.scala 39:30]
  wire  _T_84; // @[LZD.scala 39:27]
  wire  _T_85; // @[LZD.scala 39:25]
  wire  _T_87; // @[Shift.scala 12:21]
  wire [2:0] _T_89; // @[Cat.scala 29:58]
  wire [2:0] _T_90; // @[LZD.scala 55:32]
  wire [2:0] _T_91; // @[LZD.scala 55:20]
  wire [3:0] _T_92; // @[Cat.scala 29:58]
  wire [3:0] _T_93; // @[convert.scala 21:22]
  wire [8:0] _T_94; // @[convert.scala 22:36]
  wire  _T_95; // @[Shift.scala 16:24]
  wire  _T_97; // @[Shift.scala 12:21]
  wire  _T_98; // @[Shift.scala 64:52]
  wire [8:0] _T_100; // @[Cat.scala 29:58]
  wire [8:0] _T_101; // @[Shift.scala 64:27]
  wire [2:0] _T_102; // @[Shift.scala 66:70]
  wire  _T_103; // @[Shift.scala 12:21]
  wire [4:0] _T_104; // @[Shift.scala 64:52]
  wire [8:0] _T_106; // @[Cat.scala 29:58]
  wire [8:0] _T_107; // @[Shift.scala 64:27]
  wire [1:0] _T_108; // @[Shift.scala 66:70]
  wire  _T_109; // @[Shift.scala 12:21]
  wire [6:0] _T_110; // @[Shift.scala 64:52]
  wire [8:0] _T_112; // @[Cat.scala 29:58]
  wire [8:0] _T_113; // @[Shift.scala 64:27]
  wire  _T_114; // @[Shift.scala 66:70]
  wire [7:0] _T_116; // @[Shift.scala 64:52]
  wire [8:0] _T_117; // @[Cat.scala 29:58]
  wire [8:0] _T_118; // @[Shift.scala 64:27]
  wire [8:0] _T_119; // @[Shift.scala 16:10]
  wire  _T_120; // @[convert.scala 23:34]
  wire [7:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_122; // @[convert.scala 25:26]
  wire [3:0] _T_124; // @[convert.scala 25:42]
  wire  _T_127; // @[convert.scala 26:67]
  wire  _T_128; // @[convert.scala 26:51]
  wire [5:0] _T_129; // @[Cat.scala 29:58]
  wire [10:0] _T_131; // @[convert.scala 29:56]
  wire  _T_132; // @[convert.scala 29:60]
  wire  _T_133; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_136; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_145; // @[convert.scala 18:24]
  wire  _T_146; // @[convert.scala 18:40]
  wire  _T_147; // @[convert.scala 18:36]
  wire [9:0] _T_148; // @[convert.scala 19:24]
  wire [9:0] _T_149; // @[convert.scala 19:43]
  wire [9:0] _T_150; // @[convert.scala 19:39]
  wire [7:0] _T_151; // @[LZD.scala 43:32]
  wire [3:0] _T_152; // @[LZD.scala 43:32]
  wire [1:0] _T_153; // @[LZD.scala 43:32]
  wire  _T_154; // @[LZD.scala 39:14]
  wire  _T_155; // @[LZD.scala 39:21]
  wire  _T_156; // @[LZD.scala 39:30]
  wire  _T_157; // @[LZD.scala 39:27]
  wire  _T_158; // @[LZD.scala 39:25]
  wire [1:0] _T_159; // @[Cat.scala 29:58]
  wire [1:0] _T_160; // @[LZD.scala 44:32]
  wire  _T_161; // @[LZD.scala 39:14]
  wire  _T_162; // @[LZD.scala 39:21]
  wire  _T_163; // @[LZD.scala 39:30]
  wire  _T_164; // @[LZD.scala 39:27]
  wire  _T_165; // @[LZD.scala 39:25]
  wire [1:0] _T_166; // @[Cat.scala 29:58]
  wire  _T_167; // @[Shift.scala 12:21]
  wire  _T_168; // @[Shift.scala 12:21]
  wire  _T_169; // @[LZD.scala 49:16]
  wire  _T_170; // @[LZD.scala 49:27]
  wire  _T_171; // @[LZD.scala 49:25]
  wire  _T_172; // @[LZD.scala 49:47]
  wire  _T_173; // @[LZD.scala 49:59]
  wire  _T_174; // @[LZD.scala 49:35]
  wire [2:0] _T_176; // @[Cat.scala 29:58]
  wire [3:0] _T_177; // @[LZD.scala 44:32]
  wire [1:0] _T_178; // @[LZD.scala 43:32]
  wire  _T_179; // @[LZD.scala 39:14]
  wire  _T_180; // @[LZD.scala 39:21]
  wire  _T_181; // @[LZD.scala 39:30]
  wire  _T_182; // @[LZD.scala 39:27]
  wire  _T_183; // @[LZD.scala 39:25]
  wire [1:0] _T_184; // @[Cat.scala 29:58]
  wire [1:0] _T_185; // @[LZD.scala 44:32]
  wire  _T_186; // @[LZD.scala 39:14]
  wire  _T_187; // @[LZD.scala 39:21]
  wire  _T_188; // @[LZD.scala 39:30]
  wire  _T_189; // @[LZD.scala 39:27]
  wire  _T_190; // @[LZD.scala 39:25]
  wire [1:0] _T_191; // @[Cat.scala 29:58]
  wire  _T_192; // @[Shift.scala 12:21]
  wire  _T_193; // @[Shift.scala 12:21]
  wire  _T_194; // @[LZD.scala 49:16]
  wire  _T_195; // @[LZD.scala 49:27]
  wire  _T_196; // @[LZD.scala 49:25]
  wire  _T_197; // @[LZD.scala 49:47]
  wire  _T_198; // @[LZD.scala 49:59]
  wire  _T_199; // @[LZD.scala 49:35]
  wire [2:0] _T_201; // @[Cat.scala 29:58]
  wire  _T_202; // @[Shift.scala 12:21]
  wire  _T_203; // @[Shift.scala 12:21]
  wire  _T_204; // @[LZD.scala 49:16]
  wire  _T_205; // @[LZD.scala 49:27]
  wire  _T_206; // @[LZD.scala 49:25]
  wire [1:0] _T_207; // @[LZD.scala 49:47]
  wire [1:0] _T_208; // @[LZD.scala 49:59]
  wire [1:0] _T_209; // @[LZD.scala 49:35]
  wire [3:0] _T_211; // @[Cat.scala 29:58]
  wire [1:0] _T_212; // @[LZD.scala 44:32]
  wire  _T_213; // @[LZD.scala 39:14]
  wire  _T_214; // @[LZD.scala 39:21]
  wire  _T_215; // @[LZD.scala 39:30]
  wire  _T_216; // @[LZD.scala 39:27]
  wire  _T_217; // @[LZD.scala 39:25]
  wire  _T_219; // @[Shift.scala 12:21]
  wire [2:0] _T_221; // @[Cat.scala 29:58]
  wire [2:0] _T_222; // @[LZD.scala 55:32]
  wire [2:0] _T_223; // @[LZD.scala 55:20]
  wire [3:0] _T_224; // @[Cat.scala 29:58]
  wire [3:0] _T_225; // @[convert.scala 21:22]
  wire [8:0] _T_226; // @[convert.scala 22:36]
  wire  _T_227; // @[Shift.scala 16:24]
  wire  _T_229; // @[Shift.scala 12:21]
  wire  _T_230; // @[Shift.scala 64:52]
  wire [8:0] _T_232; // @[Cat.scala 29:58]
  wire [8:0] _T_233; // @[Shift.scala 64:27]
  wire [2:0] _T_234; // @[Shift.scala 66:70]
  wire  _T_235; // @[Shift.scala 12:21]
  wire [4:0] _T_236; // @[Shift.scala 64:52]
  wire [8:0] _T_238; // @[Cat.scala 29:58]
  wire [8:0] _T_239; // @[Shift.scala 64:27]
  wire [1:0] _T_240; // @[Shift.scala 66:70]
  wire  _T_241; // @[Shift.scala 12:21]
  wire [6:0] _T_242; // @[Shift.scala 64:52]
  wire [8:0] _T_244; // @[Cat.scala 29:58]
  wire [8:0] _T_245; // @[Shift.scala 64:27]
  wire  _T_246; // @[Shift.scala 66:70]
  wire [7:0] _T_248; // @[Shift.scala 64:52]
  wire [8:0] _T_249; // @[Cat.scala 29:58]
  wire [8:0] _T_250; // @[Shift.scala 64:27]
  wire [8:0] _T_251; // @[Shift.scala 16:10]
  wire  _T_252; // @[convert.scala 23:34]
  wire [7:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_254; // @[convert.scala 25:26]
  wire [3:0] _T_256; // @[convert.scala 25:42]
  wire  _T_259; // @[convert.scala 26:67]
  wire  _T_260; // @[convert.scala 26:51]
  wire [5:0] _T_261; // @[Cat.scala 29:58]
  wire [10:0] _T_263; // @[convert.scala 29:56]
  wire  _T_264; // @[convert.scala 29:60]
  wire  _T_265; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_268; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_277; // @[convert.scala 18:24]
  wire  _T_278; // @[convert.scala 18:40]
  wire  _T_279; // @[convert.scala 18:36]
  wire [9:0] _T_280; // @[convert.scala 19:24]
  wire [9:0] _T_281; // @[convert.scala 19:43]
  wire [9:0] _T_282; // @[convert.scala 19:39]
  wire [7:0] _T_283; // @[LZD.scala 43:32]
  wire [3:0] _T_284; // @[LZD.scala 43:32]
  wire [1:0] _T_285; // @[LZD.scala 43:32]
  wire  _T_286; // @[LZD.scala 39:14]
  wire  _T_287; // @[LZD.scala 39:21]
  wire  _T_288; // @[LZD.scala 39:30]
  wire  _T_289; // @[LZD.scala 39:27]
  wire  _T_290; // @[LZD.scala 39:25]
  wire [1:0] _T_291; // @[Cat.scala 29:58]
  wire [1:0] _T_292; // @[LZD.scala 44:32]
  wire  _T_293; // @[LZD.scala 39:14]
  wire  _T_294; // @[LZD.scala 39:21]
  wire  _T_295; // @[LZD.scala 39:30]
  wire  _T_296; // @[LZD.scala 39:27]
  wire  _T_297; // @[LZD.scala 39:25]
  wire [1:0] _T_298; // @[Cat.scala 29:58]
  wire  _T_299; // @[Shift.scala 12:21]
  wire  _T_300; // @[Shift.scala 12:21]
  wire  _T_301; // @[LZD.scala 49:16]
  wire  _T_302; // @[LZD.scala 49:27]
  wire  _T_303; // @[LZD.scala 49:25]
  wire  _T_304; // @[LZD.scala 49:47]
  wire  _T_305; // @[LZD.scala 49:59]
  wire  _T_306; // @[LZD.scala 49:35]
  wire [2:0] _T_308; // @[Cat.scala 29:58]
  wire [3:0] _T_309; // @[LZD.scala 44:32]
  wire [1:0] _T_310; // @[LZD.scala 43:32]
  wire  _T_311; // @[LZD.scala 39:14]
  wire  _T_312; // @[LZD.scala 39:21]
  wire  _T_313; // @[LZD.scala 39:30]
  wire  _T_314; // @[LZD.scala 39:27]
  wire  _T_315; // @[LZD.scala 39:25]
  wire [1:0] _T_316; // @[Cat.scala 29:58]
  wire [1:0] _T_317; // @[LZD.scala 44:32]
  wire  _T_318; // @[LZD.scala 39:14]
  wire  _T_319; // @[LZD.scala 39:21]
  wire  _T_320; // @[LZD.scala 39:30]
  wire  _T_321; // @[LZD.scala 39:27]
  wire  _T_322; // @[LZD.scala 39:25]
  wire [1:0] _T_323; // @[Cat.scala 29:58]
  wire  _T_324; // @[Shift.scala 12:21]
  wire  _T_325; // @[Shift.scala 12:21]
  wire  _T_326; // @[LZD.scala 49:16]
  wire  _T_327; // @[LZD.scala 49:27]
  wire  _T_328; // @[LZD.scala 49:25]
  wire  _T_329; // @[LZD.scala 49:47]
  wire  _T_330; // @[LZD.scala 49:59]
  wire  _T_331; // @[LZD.scala 49:35]
  wire [2:0] _T_333; // @[Cat.scala 29:58]
  wire  _T_334; // @[Shift.scala 12:21]
  wire  _T_335; // @[Shift.scala 12:21]
  wire  _T_336; // @[LZD.scala 49:16]
  wire  _T_337; // @[LZD.scala 49:27]
  wire  _T_338; // @[LZD.scala 49:25]
  wire [1:0] _T_339; // @[LZD.scala 49:47]
  wire [1:0] _T_340; // @[LZD.scala 49:59]
  wire [1:0] _T_341; // @[LZD.scala 49:35]
  wire [3:0] _T_343; // @[Cat.scala 29:58]
  wire [1:0] _T_344; // @[LZD.scala 44:32]
  wire  _T_345; // @[LZD.scala 39:14]
  wire  _T_346; // @[LZD.scala 39:21]
  wire  _T_347; // @[LZD.scala 39:30]
  wire  _T_348; // @[LZD.scala 39:27]
  wire  _T_349; // @[LZD.scala 39:25]
  wire  _T_351; // @[Shift.scala 12:21]
  wire [2:0] _T_353; // @[Cat.scala 29:58]
  wire [2:0] _T_354; // @[LZD.scala 55:32]
  wire [2:0] _T_355; // @[LZD.scala 55:20]
  wire [3:0] _T_356; // @[Cat.scala 29:58]
  wire [3:0] _T_357; // @[convert.scala 21:22]
  wire [8:0] _T_358; // @[convert.scala 22:36]
  wire  _T_359; // @[Shift.scala 16:24]
  wire  _T_361; // @[Shift.scala 12:21]
  wire  _T_362; // @[Shift.scala 64:52]
  wire [8:0] _T_364; // @[Cat.scala 29:58]
  wire [8:0] _T_365; // @[Shift.scala 64:27]
  wire [2:0] _T_366; // @[Shift.scala 66:70]
  wire  _T_367; // @[Shift.scala 12:21]
  wire [4:0] _T_368; // @[Shift.scala 64:52]
  wire [8:0] _T_370; // @[Cat.scala 29:58]
  wire [8:0] _T_371; // @[Shift.scala 64:27]
  wire [1:0] _T_372; // @[Shift.scala 66:70]
  wire  _T_373; // @[Shift.scala 12:21]
  wire [6:0] _T_374; // @[Shift.scala 64:52]
  wire [8:0] _T_376; // @[Cat.scala 29:58]
  wire [8:0] _T_377; // @[Shift.scala 64:27]
  wire  _T_378; // @[Shift.scala 66:70]
  wire [7:0] _T_380; // @[Shift.scala 64:52]
  wire [8:0] _T_381; // @[Cat.scala 29:58]
  wire [8:0] _T_382; // @[Shift.scala 64:27]
  wire [8:0] _T_383; // @[Shift.scala 16:10]
  wire  _T_384; // @[convert.scala 23:34]
  wire [7:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_386; // @[convert.scala 25:26]
  wire [3:0] _T_388; // @[convert.scala 25:42]
  wire  _T_391; // @[convert.scala 26:67]
  wire  _T_392; // @[convert.scala 26:51]
  wire [5:0] _T_393; // @[Cat.scala 29:58]
  wire [10:0] _T_395; // @[convert.scala 29:56]
  wire  _T_396; // @[convert.scala 29:60]
  wire  _T_397; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_400; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [5:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_408; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_409; // @[PositFMA.scala 59:34]
  wire  _T_410; // @[PositFMA.scala 59:47]
  wire  _T_411; // @[PositFMA.scala 59:45]
  wire [9:0] _T_413; // @[Cat.scala 29:58]
  wire [9:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_414; // @[PositFMA.scala 60:34]
  wire  _T_415; // @[PositFMA.scala 60:47]
  wire  _T_416; // @[PositFMA.scala 60:45]
  wire [9:0] _T_418; // @[Cat.scala 29:58]
  wire [9:0] sigB; // @[PositFMA.scala 60:76]
  wire [19:0] _T_419; // @[PositFMA.scala 61:25]
  wire [19:0] sigP; // @[PositFMA.scala 61:33]
  wire [16:0] _T_420; // @[PositFMA.scala 62:29]
  wire  _T_421; // @[PositFMA.scala 62:33]
  wire  eqTwo; // @[PositFMA.scala 62:19]
  wire  _T_422; // @[PositFMA.scala 64:29]
  wire  _T_423; // @[PositFMA.scala 64:56]
  wire  _T_424; // @[PositFMA.scala 64:51]
  wire  _T_425; // @[PositFMA.scala 64:49]
  wire  eqFour; // @[PositFMA.scala 64:76]
  wire  _T_426; // @[PositFMA.scala 66:23]
  wire  geTwo; // @[PositFMA.scala 66:43]
  wire [1:0] _T_428; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 67:38]
  wire  mulSign; // @[PositFMA.scala 68:28]
  wire [6:0] _T_429; // @[PositFMA.scala 70:30]
  wire [6:0] _GEN_12; // @[PositFMA.scala 70:44]
  wire [6:0] _T_431; // @[PositFMA.scala 70:44]
  wire [6:0] mulScale; // @[PositFMA.scala 70:44]
  wire [17:0] _T_432; // @[PositFMA.scala 73:29]
  wire [16:0] _T_433; // @[PositFMA.scala 74:29]
  wire [17:0] _T_434; // @[PositFMA.scala 74:48]
  wire [17:0] mulSigTmp; // @[PositFMA.scala 71:22]
  wire  _T_436; // @[PositFMA.scala 78:39]
  wire  _T_437; // @[PositFMA.scala 78:43]
  wire [16:0] _T_438; // @[PositFMA.scala 79:39]
  wire [18:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [18:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [7:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [6:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [5:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_464; // @[PositFMA.scala 108:29]
  wire  _T_465; // @[PositFMA.scala 108:47]
  wire  _T_466; // @[PositFMA.scala 108:45]
  wire [18:0] extAddSig; // @[Cat.scala 29:58]
  wire [6:0] _GEN_13; // @[PositFMA.scala 112:39]
  wire  mulGreater; // @[PositFMA.scala 112:39]
  wire [6:0] greaterScale; // @[PositFMA.scala 113:26]
  wire [6:0] smallerScale; // @[PositFMA.scala 114:26]
  wire [6:0] _T_470; // @[PositFMA.scala 115:36]
  wire [6:0] scaleDiff; // @[PositFMA.scala 115:36]
  wire [18:0] greaterSig; // @[PositFMA.scala 116:26]
  wire [18:0] smallerSigTmp; // @[PositFMA.scala 117:26]
  wire [6:0] _T_471; // @[PositFMA.scala 118:69]
  wire  _T_472; // @[Shift.scala 39:24]
  wire [4:0] _T_473; // @[Shift.scala 40:44]
  wire [2:0] _T_474; // @[Shift.scala 90:30]
  wire [15:0] _T_475; // @[Shift.scala 90:48]
  wire  _T_476; // @[Shift.scala 90:57]
  wire [2:0] _GEN_14; // @[Shift.scala 90:39]
  wire [2:0] _T_477; // @[Shift.scala 90:39]
  wire  _T_478; // @[Shift.scala 12:21]
  wire  _T_479; // @[Shift.scala 12:21]
  wire [15:0] _T_481; // @[Bitwise.scala 71:12]
  wire [18:0] _T_482; // @[Cat.scala 29:58]
  wire [18:0] _T_483; // @[Shift.scala 91:22]
  wire [3:0] _T_484; // @[Shift.scala 92:77]
  wire [10:0] _T_485; // @[Shift.scala 90:30]
  wire [7:0] _T_486; // @[Shift.scala 90:48]
  wire  _T_487; // @[Shift.scala 90:57]
  wire [10:0] _GEN_15; // @[Shift.scala 90:39]
  wire [10:0] _T_488; // @[Shift.scala 90:39]
  wire  _T_489; // @[Shift.scala 12:21]
  wire  _T_490; // @[Shift.scala 12:21]
  wire [7:0] _T_492; // @[Bitwise.scala 71:12]
  wire [18:0] _T_493; // @[Cat.scala 29:58]
  wire [18:0] _T_494; // @[Shift.scala 91:22]
  wire [2:0] _T_495; // @[Shift.scala 92:77]
  wire [14:0] _T_496; // @[Shift.scala 90:30]
  wire [3:0] _T_497; // @[Shift.scala 90:48]
  wire  _T_498; // @[Shift.scala 90:57]
  wire [14:0] _GEN_16; // @[Shift.scala 90:39]
  wire [14:0] _T_499; // @[Shift.scala 90:39]
  wire  _T_500; // @[Shift.scala 12:21]
  wire  _T_501; // @[Shift.scala 12:21]
  wire [3:0] _T_503; // @[Bitwise.scala 71:12]
  wire [18:0] _T_504; // @[Cat.scala 29:58]
  wire [18:0] _T_505; // @[Shift.scala 91:22]
  wire [1:0] _T_506; // @[Shift.scala 92:77]
  wire [16:0] _T_507; // @[Shift.scala 90:30]
  wire [1:0] _T_508; // @[Shift.scala 90:48]
  wire  _T_509; // @[Shift.scala 90:57]
  wire [16:0] _GEN_17; // @[Shift.scala 90:39]
  wire [16:0] _T_510; // @[Shift.scala 90:39]
  wire  _T_511; // @[Shift.scala 12:21]
  wire  _T_512; // @[Shift.scala 12:21]
  wire [1:0] _T_514; // @[Bitwise.scala 71:12]
  wire [18:0] _T_515; // @[Cat.scala 29:58]
  wire [18:0] _T_516; // @[Shift.scala 91:22]
  wire  _T_517; // @[Shift.scala 92:77]
  wire [17:0] _T_518; // @[Shift.scala 90:30]
  wire  _T_519; // @[Shift.scala 90:48]
  wire [17:0] _GEN_18; // @[Shift.scala 90:39]
  wire [17:0] _T_521; // @[Shift.scala 90:39]
  wire  _T_523; // @[Shift.scala 12:21]
  wire [18:0] _T_524; // @[Cat.scala 29:58]
  wire [18:0] _T_525; // @[Shift.scala 91:22]
  wire [18:0] _T_528; // @[Bitwise.scala 71:12]
  wire [18:0] smallerSig; // @[Shift.scala 39:10]
  wire [19:0] rawSumSig; // @[PositFMA.scala 119:34]
  wire  _T_529; // @[PositFMA.scala 120:42]
  wire  _T_530; // @[PositFMA.scala 120:46]
  wire  _T_531; // @[PositFMA.scala 120:79]
  wire  sumSign; // @[PositFMA.scala 120:63]
  wire [18:0] _T_533; // @[PositFMA.scala 121:50]
  wire [19:0] signSumSig; // @[Cat.scala 29:58]
  wire [18:0] _T_534; // @[PositFMA.scala 125:33]
  wire [18:0] _T_535; // @[PositFMA.scala 125:68]
  wire [18:0] sumXor; // @[PositFMA.scala 125:51]
  wire [15:0] _T_536; // @[LZD.scala 43:32]
  wire [7:0] _T_537; // @[LZD.scala 43:32]
  wire [3:0] _T_538; // @[LZD.scala 43:32]
  wire [1:0] _T_539; // @[LZD.scala 43:32]
  wire  _T_540; // @[LZD.scala 39:14]
  wire  _T_541; // @[LZD.scala 39:21]
  wire  _T_542; // @[LZD.scala 39:30]
  wire  _T_543; // @[LZD.scala 39:27]
  wire  _T_544; // @[LZD.scala 39:25]
  wire [1:0] _T_545; // @[Cat.scala 29:58]
  wire [1:0] _T_546; // @[LZD.scala 44:32]
  wire  _T_547; // @[LZD.scala 39:14]
  wire  _T_548; // @[LZD.scala 39:21]
  wire  _T_549; // @[LZD.scala 39:30]
  wire  _T_550; // @[LZD.scala 39:27]
  wire  _T_551; // @[LZD.scala 39:25]
  wire [1:0] _T_552; // @[Cat.scala 29:58]
  wire  _T_553; // @[Shift.scala 12:21]
  wire  _T_554; // @[Shift.scala 12:21]
  wire  _T_555; // @[LZD.scala 49:16]
  wire  _T_556; // @[LZD.scala 49:27]
  wire  _T_557; // @[LZD.scala 49:25]
  wire  _T_558; // @[LZD.scala 49:47]
  wire  _T_559; // @[LZD.scala 49:59]
  wire  _T_560; // @[LZD.scala 49:35]
  wire [2:0] _T_562; // @[Cat.scala 29:58]
  wire [3:0] _T_563; // @[LZD.scala 44:32]
  wire [1:0] _T_564; // @[LZD.scala 43:32]
  wire  _T_565; // @[LZD.scala 39:14]
  wire  _T_566; // @[LZD.scala 39:21]
  wire  _T_567; // @[LZD.scala 39:30]
  wire  _T_568; // @[LZD.scala 39:27]
  wire  _T_569; // @[LZD.scala 39:25]
  wire [1:0] _T_570; // @[Cat.scala 29:58]
  wire [1:0] _T_571; // @[LZD.scala 44:32]
  wire  _T_572; // @[LZD.scala 39:14]
  wire  _T_573; // @[LZD.scala 39:21]
  wire  _T_574; // @[LZD.scala 39:30]
  wire  _T_575; // @[LZD.scala 39:27]
  wire  _T_576; // @[LZD.scala 39:25]
  wire [1:0] _T_577; // @[Cat.scala 29:58]
  wire  _T_578; // @[Shift.scala 12:21]
  wire  _T_579; // @[Shift.scala 12:21]
  wire  _T_580; // @[LZD.scala 49:16]
  wire  _T_581; // @[LZD.scala 49:27]
  wire  _T_582; // @[LZD.scala 49:25]
  wire  _T_583; // @[LZD.scala 49:47]
  wire  _T_584; // @[LZD.scala 49:59]
  wire  _T_585; // @[LZD.scala 49:35]
  wire [2:0] _T_587; // @[Cat.scala 29:58]
  wire  _T_588; // @[Shift.scala 12:21]
  wire  _T_589; // @[Shift.scala 12:21]
  wire  _T_590; // @[LZD.scala 49:16]
  wire  _T_591; // @[LZD.scala 49:27]
  wire  _T_592; // @[LZD.scala 49:25]
  wire [1:0] _T_593; // @[LZD.scala 49:47]
  wire [1:0] _T_594; // @[LZD.scala 49:59]
  wire [1:0] _T_595; // @[LZD.scala 49:35]
  wire [3:0] _T_597; // @[Cat.scala 29:58]
  wire [7:0] _T_598; // @[LZD.scala 44:32]
  wire [3:0] _T_599; // @[LZD.scala 43:32]
  wire [1:0] _T_600; // @[LZD.scala 43:32]
  wire  _T_601; // @[LZD.scala 39:14]
  wire  _T_602; // @[LZD.scala 39:21]
  wire  _T_603; // @[LZD.scala 39:30]
  wire  _T_604; // @[LZD.scala 39:27]
  wire  _T_605; // @[LZD.scala 39:25]
  wire [1:0] _T_606; // @[Cat.scala 29:58]
  wire [1:0] _T_607; // @[LZD.scala 44:32]
  wire  _T_608; // @[LZD.scala 39:14]
  wire  _T_609; // @[LZD.scala 39:21]
  wire  _T_610; // @[LZD.scala 39:30]
  wire  _T_611; // @[LZD.scala 39:27]
  wire  _T_612; // @[LZD.scala 39:25]
  wire [1:0] _T_613; // @[Cat.scala 29:58]
  wire  _T_614; // @[Shift.scala 12:21]
  wire  _T_615; // @[Shift.scala 12:21]
  wire  _T_616; // @[LZD.scala 49:16]
  wire  _T_617; // @[LZD.scala 49:27]
  wire  _T_618; // @[LZD.scala 49:25]
  wire  _T_619; // @[LZD.scala 49:47]
  wire  _T_620; // @[LZD.scala 49:59]
  wire  _T_621; // @[LZD.scala 49:35]
  wire [2:0] _T_623; // @[Cat.scala 29:58]
  wire [3:0] _T_624; // @[LZD.scala 44:32]
  wire [1:0] _T_625; // @[LZD.scala 43:32]
  wire  _T_626; // @[LZD.scala 39:14]
  wire  _T_627; // @[LZD.scala 39:21]
  wire  _T_628; // @[LZD.scala 39:30]
  wire  _T_629; // @[LZD.scala 39:27]
  wire  _T_630; // @[LZD.scala 39:25]
  wire [1:0] _T_631; // @[Cat.scala 29:58]
  wire [1:0] _T_632; // @[LZD.scala 44:32]
  wire  _T_633; // @[LZD.scala 39:14]
  wire  _T_634; // @[LZD.scala 39:21]
  wire  _T_635; // @[LZD.scala 39:30]
  wire  _T_636; // @[LZD.scala 39:27]
  wire  _T_637; // @[LZD.scala 39:25]
  wire [1:0] _T_638; // @[Cat.scala 29:58]
  wire  _T_639; // @[Shift.scala 12:21]
  wire  _T_640; // @[Shift.scala 12:21]
  wire  _T_641; // @[LZD.scala 49:16]
  wire  _T_642; // @[LZD.scala 49:27]
  wire  _T_643; // @[LZD.scala 49:25]
  wire  _T_644; // @[LZD.scala 49:47]
  wire  _T_645; // @[LZD.scala 49:59]
  wire  _T_646; // @[LZD.scala 49:35]
  wire [2:0] _T_648; // @[Cat.scala 29:58]
  wire  _T_649; // @[Shift.scala 12:21]
  wire  _T_650; // @[Shift.scala 12:21]
  wire  _T_651; // @[LZD.scala 49:16]
  wire  _T_652; // @[LZD.scala 49:27]
  wire  _T_653; // @[LZD.scala 49:25]
  wire [1:0] _T_654; // @[LZD.scala 49:47]
  wire [1:0] _T_655; // @[LZD.scala 49:59]
  wire [1:0] _T_656; // @[LZD.scala 49:35]
  wire [3:0] _T_658; // @[Cat.scala 29:58]
  wire  _T_659; // @[Shift.scala 12:21]
  wire  _T_660; // @[Shift.scala 12:21]
  wire  _T_661; // @[LZD.scala 49:16]
  wire  _T_662; // @[LZD.scala 49:27]
  wire  _T_663; // @[LZD.scala 49:25]
  wire [2:0] _T_664; // @[LZD.scala 49:47]
  wire [2:0] _T_665; // @[LZD.scala 49:59]
  wire [2:0] _T_666; // @[LZD.scala 49:35]
  wire [4:0] _T_668; // @[Cat.scala 29:58]
  wire [2:0] _T_669; // @[LZD.scala 44:32]
  wire [1:0] _T_670; // @[LZD.scala 43:32]
  wire  _T_671; // @[LZD.scala 39:14]
  wire  _T_672; // @[LZD.scala 39:21]
  wire  _T_673; // @[LZD.scala 39:30]
  wire  _T_674; // @[LZD.scala 39:27]
  wire  _T_675; // @[LZD.scala 39:25]
  wire [1:0] _T_676; // @[Cat.scala 29:58]
  wire  _T_677; // @[LZD.scala 44:32]
  wire  _T_679; // @[Shift.scala 12:21]
  wire  _T_681; // @[LZD.scala 55:32]
  wire  _T_682; // @[LZD.scala 55:20]
  wire  _T_684; // @[Shift.scala 12:21]
  wire [3:0] _T_687; // @[Cat.scala 29:58]
  wire [3:0] _T_688; // @[LZD.scala 55:32]
  wire [3:0] _T_689; // @[LZD.scala 55:20]
  wire [4:0] sumLZD; // @[Cat.scala 29:58]
  wire [4:0] shiftValue; // @[PositFMA.scala 127:24]
  wire [17:0] _T_690; // @[PositFMA.scala 128:38]
  wire  _T_691; // @[Shift.scala 16:24]
  wire  _T_693; // @[Shift.scala 12:21]
  wire [1:0] _T_694; // @[Shift.scala 64:52]
  wire [17:0] _T_696; // @[Cat.scala 29:58]
  wire [17:0] _T_697; // @[Shift.scala 64:27]
  wire [3:0] _T_698; // @[Shift.scala 66:70]
  wire  _T_699; // @[Shift.scala 12:21]
  wire [9:0] _T_700; // @[Shift.scala 64:52]
  wire [17:0] _T_702; // @[Cat.scala 29:58]
  wire [17:0] _T_703; // @[Shift.scala 64:27]
  wire [2:0] _T_704; // @[Shift.scala 66:70]
  wire  _T_705; // @[Shift.scala 12:21]
  wire [13:0] _T_706; // @[Shift.scala 64:52]
  wire [17:0] _T_708; // @[Cat.scala 29:58]
  wire [17:0] _T_709; // @[Shift.scala 64:27]
  wire [1:0] _T_710; // @[Shift.scala 66:70]
  wire  _T_711; // @[Shift.scala 12:21]
  wire [15:0] _T_712; // @[Shift.scala 64:52]
  wire [17:0] _T_714; // @[Cat.scala 29:58]
  wire [17:0] _T_715; // @[Shift.scala 64:27]
  wire  _T_716; // @[Shift.scala 66:70]
  wire [16:0] _T_718; // @[Shift.scala 64:52]
  wire [17:0] _T_719; // @[Cat.scala 29:58]
  wire [17:0] _T_720; // @[Shift.scala 64:27]
  wire [17:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [6:0] _T_722; // @[PositFMA.scala 131:36]
  wire [6:0] _T_723; // @[PositFMA.scala 131:36]
  wire [5:0] _T_724; // @[Cat.scala 29:58]
  wire [5:0] _T_725; // @[PositFMA.scala 131:61]
  wire [6:0] _GEN_19; // @[PositFMA.scala 131:42]
  wire [6:0] _T_727; // @[PositFMA.scala 131:42]
  wire [6:0] sumScale; // @[PositFMA.scala 131:42]
  wire [7:0] sumFrac; // @[PositFMA.scala 132:41]
  wire [9:0] grsTmp; // @[PositFMA.scala 135:41]
  wire [1:0] _T_728; // @[PositFMA.scala 138:40]
  wire [7:0] _T_729; // @[PositFMA.scala 138:56]
  wire  _T_730; // @[PositFMA.scala 138:60]
  wire  underflow; // @[PositFMA.scala 145:32]
  wire  overflow; // @[PositFMA.scala 146:32]
  wire  _T_731; // @[PositFMA.scala 155:32]
  wire  decF_isZero; // @[PositFMA.scala 155:20]
  wire [6:0] _T_733; // @[Mux.scala 87:16]
  wire [6:0] _T_734; // @[Mux.scala 87:16]
  wire [5:0] _GEN_20; // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  wire [5:0] decF_scale; // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  wire  _T_735; // @[convert.scala 46:61]
  wire  _T_736; // @[convert.scala 46:52]
  wire  _T_738; // @[convert.scala 46:42]
  wire [4:0] _T_739; // @[convert.scala 48:34]
  wire  _T_740; // @[convert.scala 49:36]
  wire [4:0] _T_742; // @[convert.scala 50:36]
  wire [4:0] _T_743; // @[convert.scala 50:36]
  wire [4:0] _T_744; // @[convert.scala 50:28]
  wire  _T_745; // @[convert.scala 51:31]
  wire  _T_746; // @[convert.scala 52:43]
  wire [13:0] _T_750; // @[Cat.scala 29:58]
  wire [4:0] _T_751; // @[Shift.scala 39:17]
  wire  _T_752; // @[Shift.scala 39:24]
  wire [3:0] _T_753; // @[Shift.scala 40:44]
  wire [5:0] _T_754; // @[Shift.scala 90:30]
  wire [7:0] _T_755; // @[Shift.scala 90:48]
  wire  _T_756; // @[Shift.scala 90:57]
  wire [5:0] _GEN_21; // @[Shift.scala 90:39]
  wire [5:0] _T_757; // @[Shift.scala 90:39]
  wire  _T_758; // @[Shift.scala 12:21]
  wire  _T_759; // @[Shift.scala 12:21]
  wire [7:0] _T_761; // @[Bitwise.scala 71:12]
  wire [13:0] _T_762; // @[Cat.scala 29:58]
  wire [13:0] _T_763; // @[Shift.scala 91:22]
  wire [2:0] _T_764; // @[Shift.scala 92:77]
  wire [9:0] _T_765; // @[Shift.scala 90:30]
  wire [3:0] _T_766; // @[Shift.scala 90:48]
  wire  _T_767; // @[Shift.scala 90:57]
  wire [9:0] _GEN_22; // @[Shift.scala 90:39]
  wire [9:0] _T_768; // @[Shift.scala 90:39]
  wire  _T_769; // @[Shift.scala 12:21]
  wire  _T_770; // @[Shift.scala 12:21]
  wire [3:0] _T_772; // @[Bitwise.scala 71:12]
  wire [13:0] _T_773; // @[Cat.scala 29:58]
  wire [13:0] _T_774; // @[Shift.scala 91:22]
  wire [1:0] _T_775; // @[Shift.scala 92:77]
  wire [11:0] _T_776; // @[Shift.scala 90:30]
  wire [1:0] _T_777; // @[Shift.scala 90:48]
  wire  _T_778; // @[Shift.scala 90:57]
  wire [11:0] _GEN_23; // @[Shift.scala 90:39]
  wire [11:0] _T_779; // @[Shift.scala 90:39]
  wire  _T_780; // @[Shift.scala 12:21]
  wire  _T_781; // @[Shift.scala 12:21]
  wire [1:0] _T_783; // @[Bitwise.scala 71:12]
  wire [13:0] _T_784; // @[Cat.scala 29:58]
  wire [13:0] _T_785; // @[Shift.scala 91:22]
  wire  _T_786; // @[Shift.scala 92:77]
  wire [12:0] _T_787; // @[Shift.scala 90:30]
  wire  _T_788; // @[Shift.scala 90:48]
  wire [12:0] _GEN_24; // @[Shift.scala 90:39]
  wire [12:0] _T_790; // @[Shift.scala 90:39]
  wire  _T_792; // @[Shift.scala 12:21]
  wire [13:0] _T_793; // @[Cat.scala 29:58]
  wire [13:0] _T_794; // @[Shift.scala 91:22]
  wire [13:0] _T_797; // @[Bitwise.scala 71:12]
  wire [13:0] _T_798; // @[Shift.scala 39:10]
  wire  _T_799; // @[convert.scala 55:31]
  wire  _T_800; // @[convert.scala 56:31]
  wire  _T_801; // @[convert.scala 57:31]
  wire  _T_802; // @[convert.scala 58:31]
  wire [10:0] _T_803; // @[convert.scala 59:69]
  wire  _T_804; // @[convert.scala 59:81]
  wire  _T_805; // @[convert.scala 59:50]
  wire  _T_807; // @[convert.scala 60:81]
  wire  _T_808; // @[convert.scala 61:44]
  wire  _T_809; // @[convert.scala 61:52]
  wire  _T_810; // @[convert.scala 61:36]
  wire  _T_811; // @[convert.scala 62:63]
  wire  _T_812; // @[convert.scala 62:103]
  wire  _T_813; // @[convert.scala 62:60]
  wire [10:0] _GEN_25; // @[convert.scala 63:56]
  wire [10:0] _T_816; // @[convert.scala 63:56]
  wire [11:0] _T_817; // @[Cat.scala 29:58]
  reg  _T_821; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [11:0] _T_825; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 12'hfff : 12'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{11'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 12'hfff : 12'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{11'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[11]; // @[convert.scala 18:24]
  assign _T_14 = realA[10]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[10:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[9:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[9:2]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[7:4]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20[3:2]; // @[LZD.scala 43:32]
  assign _T_22 = _T_21 != 2'h0; // @[LZD.scala 39:14]
  assign _T_23 = _T_21[1]; // @[LZD.scala 39:21]
  assign _T_24 = _T_21[0]; // @[LZD.scala 39:30]
  assign _T_25 = ~ _T_24; // @[LZD.scala 39:27]
  assign _T_26 = _T_23 | _T_25; // @[LZD.scala 39:25]
  assign _T_27 = {_T_22,_T_26}; // @[Cat.scala 29:58]
  assign _T_28 = _T_20[1:0]; // @[LZD.scala 44:32]
  assign _T_29 = _T_28 != 2'h0; // @[LZD.scala 39:14]
  assign _T_30 = _T_28[1]; // @[LZD.scala 39:21]
  assign _T_31 = _T_28[0]; // @[LZD.scala 39:30]
  assign _T_32 = ~ _T_31; // @[LZD.scala 39:27]
  assign _T_33 = _T_30 | _T_32; // @[LZD.scala 39:25]
  assign _T_34 = {_T_29,_T_33}; // @[Cat.scala 29:58]
  assign _T_35 = _T_27[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_34[1]; // @[Shift.scala 12:21]
  assign _T_37 = _T_35 | _T_36; // @[LZD.scala 49:16]
  assign _T_38 = ~ _T_36; // @[LZD.scala 49:27]
  assign _T_39 = _T_35 | _T_38; // @[LZD.scala 49:25]
  assign _T_40 = _T_27[0:0]; // @[LZD.scala 49:47]
  assign _T_41 = _T_34[0:0]; // @[LZD.scala 49:59]
  assign _T_42 = _T_35 ? _T_40 : _T_41; // @[LZD.scala 49:35]
  assign _T_44 = {_T_37,_T_39,_T_42}; // @[Cat.scala 29:58]
  assign _T_45 = _T_19[3:0]; // @[LZD.scala 44:32]
  assign _T_46 = _T_45[3:2]; // @[LZD.scala 43:32]
  assign _T_47 = _T_46 != 2'h0; // @[LZD.scala 39:14]
  assign _T_48 = _T_46[1]; // @[LZD.scala 39:21]
  assign _T_49 = _T_46[0]; // @[LZD.scala 39:30]
  assign _T_50 = ~ _T_49; // @[LZD.scala 39:27]
  assign _T_51 = _T_48 | _T_50; // @[LZD.scala 39:25]
  assign _T_52 = {_T_47,_T_51}; // @[Cat.scala 29:58]
  assign _T_53 = _T_45[1:0]; // @[LZD.scala 44:32]
  assign _T_54 = _T_53 != 2'h0; // @[LZD.scala 39:14]
  assign _T_55 = _T_53[1]; // @[LZD.scala 39:21]
  assign _T_56 = _T_53[0]; // @[LZD.scala 39:30]
  assign _T_57 = ~ _T_56; // @[LZD.scala 39:27]
  assign _T_58 = _T_55 | _T_57; // @[LZD.scala 39:25]
  assign _T_59 = {_T_54,_T_58}; // @[Cat.scala 29:58]
  assign _T_60 = _T_52[1]; // @[Shift.scala 12:21]
  assign _T_61 = _T_59[1]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60 | _T_61; // @[LZD.scala 49:16]
  assign _T_63 = ~ _T_61; // @[LZD.scala 49:27]
  assign _T_64 = _T_60 | _T_63; // @[LZD.scala 49:25]
  assign _T_65 = _T_52[0:0]; // @[LZD.scala 49:47]
  assign _T_66 = _T_59[0:0]; // @[LZD.scala 49:59]
  assign _T_67 = _T_60 ? _T_65 : _T_66; // @[LZD.scala 49:35]
  assign _T_69 = {_T_62,_T_64,_T_67}; // @[Cat.scala 29:58]
  assign _T_70 = _T_44[2]; // @[Shift.scala 12:21]
  assign _T_71 = _T_69[2]; // @[Shift.scala 12:21]
  assign _T_72 = _T_70 | _T_71; // @[LZD.scala 49:16]
  assign _T_73 = ~ _T_71; // @[LZD.scala 49:27]
  assign _T_74 = _T_70 | _T_73; // @[LZD.scala 49:25]
  assign _T_75 = _T_44[1:0]; // @[LZD.scala 49:47]
  assign _T_76 = _T_69[1:0]; // @[LZD.scala 49:59]
  assign _T_77 = _T_70 ? _T_75 : _T_76; // @[LZD.scala 49:35]
  assign _T_79 = {_T_72,_T_74,_T_77}; // @[Cat.scala 29:58]
  assign _T_80 = _T_18[1:0]; // @[LZD.scala 44:32]
  assign _T_81 = _T_80 != 2'h0; // @[LZD.scala 39:14]
  assign _T_82 = _T_80[1]; // @[LZD.scala 39:21]
  assign _T_83 = _T_80[0]; // @[LZD.scala 39:30]
  assign _T_84 = ~ _T_83; // @[LZD.scala 39:27]
  assign _T_85 = _T_82 | _T_84; // @[LZD.scala 39:25]
  assign _T_87 = _T_79[3]; // @[Shift.scala 12:21]
  assign _T_89 = {1'h1,_T_81,_T_85}; // @[Cat.scala 29:58]
  assign _T_90 = _T_79[2:0]; // @[LZD.scala 55:32]
  assign _T_91 = _T_87 ? _T_90 : _T_89; // @[LZD.scala 55:20]
  assign _T_92 = {_T_87,_T_91}; // @[Cat.scala 29:58]
  assign _T_93 = ~ _T_92; // @[convert.scala 21:22]
  assign _T_94 = realA[8:0]; // @[convert.scala 22:36]
  assign _T_95 = _T_93 < 4'h9; // @[Shift.scala 16:24]
  assign _T_97 = _T_93[3]; // @[Shift.scala 12:21]
  assign _T_98 = _T_94[0:0]; // @[Shift.scala 64:52]
  assign _T_100 = {_T_98,8'h0}; // @[Cat.scala 29:58]
  assign _T_101 = _T_97 ? _T_100 : _T_94; // @[Shift.scala 64:27]
  assign _T_102 = _T_93[2:0]; // @[Shift.scala 66:70]
  assign _T_103 = _T_102[2]; // @[Shift.scala 12:21]
  assign _T_104 = _T_101[4:0]; // @[Shift.scala 64:52]
  assign _T_106 = {_T_104,4'h0}; // @[Cat.scala 29:58]
  assign _T_107 = _T_103 ? _T_106 : _T_101; // @[Shift.scala 64:27]
  assign _T_108 = _T_102[1:0]; // @[Shift.scala 66:70]
  assign _T_109 = _T_108[1]; // @[Shift.scala 12:21]
  assign _T_110 = _T_107[6:0]; // @[Shift.scala 64:52]
  assign _T_112 = {_T_110,2'h0}; // @[Cat.scala 29:58]
  assign _T_113 = _T_109 ? _T_112 : _T_107; // @[Shift.scala 64:27]
  assign _T_114 = _T_108[0:0]; // @[Shift.scala 66:70]
  assign _T_116 = _T_113[7:0]; // @[Shift.scala 64:52]
  assign _T_117 = {_T_116,1'h0}; // @[Cat.scala 29:58]
  assign _T_118 = _T_114 ? _T_117 : _T_113; // @[Shift.scala 64:27]
  assign _T_119 = _T_95 ? _T_118 : 9'h0; // @[Shift.scala 16:10]
  assign _T_120 = _T_119[8:8]; // @[convert.scala 23:34]
  assign decA_fraction = _T_119[7:0]; // @[convert.scala 24:34]
  assign _T_122 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_124 = _T_15 ? _T_93 : _T_92; // @[convert.scala 25:42]
  assign _T_127 = ~ _T_120; // @[convert.scala 26:67]
  assign _T_128 = _T_13 ? _T_127 : _T_120; // @[convert.scala 26:51]
  assign _T_129 = {_T_122,_T_124,_T_128}; // @[Cat.scala 29:58]
  assign _T_131 = realA[10:0]; // @[convert.scala 29:56]
  assign _T_132 = _T_131 != 11'h0; // @[convert.scala 29:60]
  assign _T_133 = ~ _T_132; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_133; // @[convert.scala 29:39]
  assign _T_136 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_136 & _T_133; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_129); // @[convert.scala 32:24]
  assign _T_145 = io_B[11]; // @[convert.scala 18:24]
  assign _T_146 = io_B[10]; // @[convert.scala 18:40]
  assign _T_147 = _T_145 ^ _T_146; // @[convert.scala 18:36]
  assign _T_148 = io_B[10:1]; // @[convert.scala 19:24]
  assign _T_149 = io_B[9:0]; // @[convert.scala 19:43]
  assign _T_150 = _T_148 ^ _T_149; // @[convert.scala 19:39]
  assign _T_151 = _T_150[9:2]; // @[LZD.scala 43:32]
  assign _T_152 = _T_151[7:4]; // @[LZD.scala 43:32]
  assign _T_153 = _T_152[3:2]; // @[LZD.scala 43:32]
  assign _T_154 = _T_153 != 2'h0; // @[LZD.scala 39:14]
  assign _T_155 = _T_153[1]; // @[LZD.scala 39:21]
  assign _T_156 = _T_153[0]; // @[LZD.scala 39:30]
  assign _T_157 = ~ _T_156; // @[LZD.scala 39:27]
  assign _T_158 = _T_155 | _T_157; // @[LZD.scala 39:25]
  assign _T_159 = {_T_154,_T_158}; // @[Cat.scala 29:58]
  assign _T_160 = _T_152[1:0]; // @[LZD.scala 44:32]
  assign _T_161 = _T_160 != 2'h0; // @[LZD.scala 39:14]
  assign _T_162 = _T_160[1]; // @[LZD.scala 39:21]
  assign _T_163 = _T_160[0]; // @[LZD.scala 39:30]
  assign _T_164 = ~ _T_163; // @[LZD.scala 39:27]
  assign _T_165 = _T_162 | _T_164; // @[LZD.scala 39:25]
  assign _T_166 = {_T_161,_T_165}; // @[Cat.scala 29:58]
  assign _T_167 = _T_159[1]; // @[Shift.scala 12:21]
  assign _T_168 = _T_166[1]; // @[Shift.scala 12:21]
  assign _T_169 = _T_167 | _T_168; // @[LZD.scala 49:16]
  assign _T_170 = ~ _T_168; // @[LZD.scala 49:27]
  assign _T_171 = _T_167 | _T_170; // @[LZD.scala 49:25]
  assign _T_172 = _T_159[0:0]; // @[LZD.scala 49:47]
  assign _T_173 = _T_166[0:0]; // @[LZD.scala 49:59]
  assign _T_174 = _T_167 ? _T_172 : _T_173; // @[LZD.scala 49:35]
  assign _T_176 = {_T_169,_T_171,_T_174}; // @[Cat.scala 29:58]
  assign _T_177 = _T_151[3:0]; // @[LZD.scala 44:32]
  assign _T_178 = _T_177[3:2]; // @[LZD.scala 43:32]
  assign _T_179 = _T_178 != 2'h0; // @[LZD.scala 39:14]
  assign _T_180 = _T_178[1]; // @[LZD.scala 39:21]
  assign _T_181 = _T_178[0]; // @[LZD.scala 39:30]
  assign _T_182 = ~ _T_181; // @[LZD.scala 39:27]
  assign _T_183 = _T_180 | _T_182; // @[LZD.scala 39:25]
  assign _T_184 = {_T_179,_T_183}; // @[Cat.scala 29:58]
  assign _T_185 = _T_177[1:0]; // @[LZD.scala 44:32]
  assign _T_186 = _T_185 != 2'h0; // @[LZD.scala 39:14]
  assign _T_187 = _T_185[1]; // @[LZD.scala 39:21]
  assign _T_188 = _T_185[0]; // @[LZD.scala 39:30]
  assign _T_189 = ~ _T_188; // @[LZD.scala 39:27]
  assign _T_190 = _T_187 | _T_189; // @[LZD.scala 39:25]
  assign _T_191 = {_T_186,_T_190}; // @[Cat.scala 29:58]
  assign _T_192 = _T_184[1]; // @[Shift.scala 12:21]
  assign _T_193 = _T_191[1]; // @[Shift.scala 12:21]
  assign _T_194 = _T_192 | _T_193; // @[LZD.scala 49:16]
  assign _T_195 = ~ _T_193; // @[LZD.scala 49:27]
  assign _T_196 = _T_192 | _T_195; // @[LZD.scala 49:25]
  assign _T_197 = _T_184[0:0]; // @[LZD.scala 49:47]
  assign _T_198 = _T_191[0:0]; // @[LZD.scala 49:59]
  assign _T_199 = _T_192 ? _T_197 : _T_198; // @[LZD.scala 49:35]
  assign _T_201 = {_T_194,_T_196,_T_199}; // @[Cat.scala 29:58]
  assign _T_202 = _T_176[2]; // @[Shift.scala 12:21]
  assign _T_203 = _T_201[2]; // @[Shift.scala 12:21]
  assign _T_204 = _T_202 | _T_203; // @[LZD.scala 49:16]
  assign _T_205 = ~ _T_203; // @[LZD.scala 49:27]
  assign _T_206 = _T_202 | _T_205; // @[LZD.scala 49:25]
  assign _T_207 = _T_176[1:0]; // @[LZD.scala 49:47]
  assign _T_208 = _T_201[1:0]; // @[LZD.scala 49:59]
  assign _T_209 = _T_202 ? _T_207 : _T_208; // @[LZD.scala 49:35]
  assign _T_211 = {_T_204,_T_206,_T_209}; // @[Cat.scala 29:58]
  assign _T_212 = _T_150[1:0]; // @[LZD.scala 44:32]
  assign _T_213 = _T_212 != 2'h0; // @[LZD.scala 39:14]
  assign _T_214 = _T_212[1]; // @[LZD.scala 39:21]
  assign _T_215 = _T_212[0]; // @[LZD.scala 39:30]
  assign _T_216 = ~ _T_215; // @[LZD.scala 39:27]
  assign _T_217 = _T_214 | _T_216; // @[LZD.scala 39:25]
  assign _T_219 = _T_211[3]; // @[Shift.scala 12:21]
  assign _T_221 = {1'h1,_T_213,_T_217}; // @[Cat.scala 29:58]
  assign _T_222 = _T_211[2:0]; // @[LZD.scala 55:32]
  assign _T_223 = _T_219 ? _T_222 : _T_221; // @[LZD.scala 55:20]
  assign _T_224 = {_T_219,_T_223}; // @[Cat.scala 29:58]
  assign _T_225 = ~ _T_224; // @[convert.scala 21:22]
  assign _T_226 = io_B[8:0]; // @[convert.scala 22:36]
  assign _T_227 = _T_225 < 4'h9; // @[Shift.scala 16:24]
  assign _T_229 = _T_225[3]; // @[Shift.scala 12:21]
  assign _T_230 = _T_226[0:0]; // @[Shift.scala 64:52]
  assign _T_232 = {_T_230,8'h0}; // @[Cat.scala 29:58]
  assign _T_233 = _T_229 ? _T_232 : _T_226; // @[Shift.scala 64:27]
  assign _T_234 = _T_225[2:0]; // @[Shift.scala 66:70]
  assign _T_235 = _T_234[2]; // @[Shift.scala 12:21]
  assign _T_236 = _T_233[4:0]; // @[Shift.scala 64:52]
  assign _T_238 = {_T_236,4'h0}; // @[Cat.scala 29:58]
  assign _T_239 = _T_235 ? _T_238 : _T_233; // @[Shift.scala 64:27]
  assign _T_240 = _T_234[1:0]; // @[Shift.scala 66:70]
  assign _T_241 = _T_240[1]; // @[Shift.scala 12:21]
  assign _T_242 = _T_239[6:0]; // @[Shift.scala 64:52]
  assign _T_244 = {_T_242,2'h0}; // @[Cat.scala 29:58]
  assign _T_245 = _T_241 ? _T_244 : _T_239; // @[Shift.scala 64:27]
  assign _T_246 = _T_240[0:0]; // @[Shift.scala 66:70]
  assign _T_248 = _T_245[7:0]; // @[Shift.scala 64:52]
  assign _T_249 = {_T_248,1'h0}; // @[Cat.scala 29:58]
  assign _T_250 = _T_246 ? _T_249 : _T_245; // @[Shift.scala 64:27]
  assign _T_251 = _T_227 ? _T_250 : 9'h0; // @[Shift.scala 16:10]
  assign _T_252 = _T_251[8:8]; // @[convert.scala 23:34]
  assign decB_fraction = _T_251[7:0]; // @[convert.scala 24:34]
  assign _T_254 = _T_147 == 1'h0; // @[convert.scala 25:26]
  assign _T_256 = _T_147 ? _T_225 : _T_224; // @[convert.scala 25:42]
  assign _T_259 = ~ _T_252; // @[convert.scala 26:67]
  assign _T_260 = _T_145 ? _T_259 : _T_252; // @[convert.scala 26:51]
  assign _T_261 = {_T_254,_T_256,_T_260}; // @[Cat.scala 29:58]
  assign _T_263 = io_B[10:0]; // @[convert.scala 29:56]
  assign _T_264 = _T_263 != 11'h0; // @[convert.scala 29:60]
  assign _T_265 = ~ _T_264; // @[convert.scala 29:41]
  assign decB_isNaR = _T_145 & _T_265; // @[convert.scala 29:39]
  assign _T_268 = _T_145 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_268 & _T_265; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_261); // @[convert.scala 32:24]
  assign _T_277 = realC[11]; // @[convert.scala 18:24]
  assign _T_278 = realC[10]; // @[convert.scala 18:40]
  assign _T_279 = _T_277 ^ _T_278; // @[convert.scala 18:36]
  assign _T_280 = realC[10:1]; // @[convert.scala 19:24]
  assign _T_281 = realC[9:0]; // @[convert.scala 19:43]
  assign _T_282 = _T_280 ^ _T_281; // @[convert.scala 19:39]
  assign _T_283 = _T_282[9:2]; // @[LZD.scala 43:32]
  assign _T_284 = _T_283[7:4]; // @[LZD.scala 43:32]
  assign _T_285 = _T_284[3:2]; // @[LZD.scala 43:32]
  assign _T_286 = _T_285 != 2'h0; // @[LZD.scala 39:14]
  assign _T_287 = _T_285[1]; // @[LZD.scala 39:21]
  assign _T_288 = _T_285[0]; // @[LZD.scala 39:30]
  assign _T_289 = ~ _T_288; // @[LZD.scala 39:27]
  assign _T_290 = _T_287 | _T_289; // @[LZD.scala 39:25]
  assign _T_291 = {_T_286,_T_290}; // @[Cat.scala 29:58]
  assign _T_292 = _T_284[1:0]; // @[LZD.scala 44:32]
  assign _T_293 = _T_292 != 2'h0; // @[LZD.scala 39:14]
  assign _T_294 = _T_292[1]; // @[LZD.scala 39:21]
  assign _T_295 = _T_292[0]; // @[LZD.scala 39:30]
  assign _T_296 = ~ _T_295; // @[LZD.scala 39:27]
  assign _T_297 = _T_294 | _T_296; // @[LZD.scala 39:25]
  assign _T_298 = {_T_293,_T_297}; // @[Cat.scala 29:58]
  assign _T_299 = _T_291[1]; // @[Shift.scala 12:21]
  assign _T_300 = _T_298[1]; // @[Shift.scala 12:21]
  assign _T_301 = _T_299 | _T_300; // @[LZD.scala 49:16]
  assign _T_302 = ~ _T_300; // @[LZD.scala 49:27]
  assign _T_303 = _T_299 | _T_302; // @[LZD.scala 49:25]
  assign _T_304 = _T_291[0:0]; // @[LZD.scala 49:47]
  assign _T_305 = _T_298[0:0]; // @[LZD.scala 49:59]
  assign _T_306 = _T_299 ? _T_304 : _T_305; // @[LZD.scala 49:35]
  assign _T_308 = {_T_301,_T_303,_T_306}; // @[Cat.scala 29:58]
  assign _T_309 = _T_283[3:0]; // @[LZD.scala 44:32]
  assign _T_310 = _T_309[3:2]; // @[LZD.scala 43:32]
  assign _T_311 = _T_310 != 2'h0; // @[LZD.scala 39:14]
  assign _T_312 = _T_310[1]; // @[LZD.scala 39:21]
  assign _T_313 = _T_310[0]; // @[LZD.scala 39:30]
  assign _T_314 = ~ _T_313; // @[LZD.scala 39:27]
  assign _T_315 = _T_312 | _T_314; // @[LZD.scala 39:25]
  assign _T_316 = {_T_311,_T_315}; // @[Cat.scala 29:58]
  assign _T_317 = _T_309[1:0]; // @[LZD.scala 44:32]
  assign _T_318 = _T_317 != 2'h0; // @[LZD.scala 39:14]
  assign _T_319 = _T_317[1]; // @[LZD.scala 39:21]
  assign _T_320 = _T_317[0]; // @[LZD.scala 39:30]
  assign _T_321 = ~ _T_320; // @[LZD.scala 39:27]
  assign _T_322 = _T_319 | _T_321; // @[LZD.scala 39:25]
  assign _T_323 = {_T_318,_T_322}; // @[Cat.scala 29:58]
  assign _T_324 = _T_316[1]; // @[Shift.scala 12:21]
  assign _T_325 = _T_323[1]; // @[Shift.scala 12:21]
  assign _T_326 = _T_324 | _T_325; // @[LZD.scala 49:16]
  assign _T_327 = ~ _T_325; // @[LZD.scala 49:27]
  assign _T_328 = _T_324 | _T_327; // @[LZD.scala 49:25]
  assign _T_329 = _T_316[0:0]; // @[LZD.scala 49:47]
  assign _T_330 = _T_323[0:0]; // @[LZD.scala 49:59]
  assign _T_331 = _T_324 ? _T_329 : _T_330; // @[LZD.scala 49:35]
  assign _T_333 = {_T_326,_T_328,_T_331}; // @[Cat.scala 29:58]
  assign _T_334 = _T_308[2]; // @[Shift.scala 12:21]
  assign _T_335 = _T_333[2]; // @[Shift.scala 12:21]
  assign _T_336 = _T_334 | _T_335; // @[LZD.scala 49:16]
  assign _T_337 = ~ _T_335; // @[LZD.scala 49:27]
  assign _T_338 = _T_334 | _T_337; // @[LZD.scala 49:25]
  assign _T_339 = _T_308[1:0]; // @[LZD.scala 49:47]
  assign _T_340 = _T_333[1:0]; // @[LZD.scala 49:59]
  assign _T_341 = _T_334 ? _T_339 : _T_340; // @[LZD.scala 49:35]
  assign _T_343 = {_T_336,_T_338,_T_341}; // @[Cat.scala 29:58]
  assign _T_344 = _T_282[1:0]; // @[LZD.scala 44:32]
  assign _T_345 = _T_344 != 2'h0; // @[LZD.scala 39:14]
  assign _T_346 = _T_344[1]; // @[LZD.scala 39:21]
  assign _T_347 = _T_344[0]; // @[LZD.scala 39:30]
  assign _T_348 = ~ _T_347; // @[LZD.scala 39:27]
  assign _T_349 = _T_346 | _T_348; // @[LZD.scala 39:25]
  assign _T_351 = _T_343[3]; // @[Shift.scala 12:21]
  assign _T_353 = {1'h1,_T_345,_T_349}; // @[Cat.scala 29:58]
  assign _T_354 = _T_343[2:0]; // @[LZD.scala 55:32]
  assign _T_355 = _T_351 ? _T_354 : _T_353; // @[LZD.scala 55:20]
  assign _T_356 = {_T_351,_T_355}; // @[Cat.scala 29:58]
  assign _T_357 = ~ _T_356; // @[convert.scala 21:22]
  assign _T_358 = realC[8:0]; // @[convert.scala 22:36]
  assign _T_359 = _T_357 < 4'h9; // @[Shift.scala 16:24]
  assign _T_361 = _T_357[3]; // @[Shift.scala 12:21]
  assign _T_362 = _T_358[0:0]; // @[Shift.scala 64:52]
  assign _T_364 = {_T_362,8'h0}; // @[Cat.scala 29:58]
  assign _T_365 = _T_361 ? _T_364 : _T_358; // @[Shift.scala 64:27]
  assign _T_366 = _T_357[2:0]; // @[Shift.scala 66:70]
  assign _T_367 = _T_366[2]; // @[Shift.scala 12:21]
  assign _T_368 = _T_365[4:0]; // @[Shift.scala 64:52]
  assign _T_370 = {_T_368,4'h0}; // @[Cat.scala 29:58]
  assign _T_371 = _T_367 ? _T_370 : _T_365; // @[Shift.scala 64:27]
  assign _T_372 = _T_366[1:0]; // @[Shift.scala 66:70]
  assign _T_373 = _T_372[1]; // @[Shift.scala 12:21]
  assign _T_374 = _T_371[6:0]; // @[Shift.scala 64:52]
  assign _T_376 = {_T_374,2'h0}; // @[Cat.scala 29:58]
  assign _T_377 = _T_373 ? _T_376 : _T_371; // @[Shift.scala 64:27]
  assign _T_378 = _T_372[0:0]; // @[Shift.scala 66:70]
  assign _T_380 = _T_377[7:0]; // @[Shift.scala 64:52]
  assign _T_381 = {_T_380,1'h0}; // @[Cat.scala 29:58]
  assign _T_382 = _T_378 ? _T_381 : _T_377; // @[Shift.scala 64:27]
  assign _T_383 = _T_359 ? _T_382 : 9'h0; // @[Shift.scala 16:10]
  assign _T_384 = _T_383[8:8]; // @[convert.scala 23:34]
  assign decC_fraction = _T_383[7:0]; // @[convert.scala 24:34]
  assign _T_386 = _T_279 == 1'h0; // @[convert.scala 25:26]
  assign _T_388 = _T_279 ? _T_357 : _T_356; // @[convert.scala 25:42]
  assign _T_391 = ~ _T_384; // @[convert.scala 26:67]
  assign _T_392 = _T_277 ? _T_391 : _T_384; // @[convert.scala 26:51]
  assign _T_393 = {_T_386,_T_388,_T_392}; // @[Cat.scala 29:58]
  assign _T_395 = realC[10:0]; // @[convert.scala 29:56]
  assign _T_396 = _T_395 != 11'h0; // @[convert.scala 29:60]
  assign _T_397 = ~ _T_396; // @[convert.scala 29:41]
  assign decC_isNaR = _T_277 & _T_397; // @[convert.scala 29:39]
  assign _T_400 = _T_277 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_400 & _T_397; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_393); // @[convert.scala 32:24]
  assign _T_408 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_408 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_409 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_410 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_411 = _T_409 & _T_410; // @[PositFMA.scala 59:45]
  assign _T_413 = {_T_13,_T_411,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_413); // @[PositFMA.scala 59:76]
  assign _T_414 = ~ _T_145; // @[PositFMA.scala 60:34]
  assign _T_415 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_416 = _T_414 & _T_415; // @[PositFMA.scala 60:45]
  assign _T_418 = {_T_145,_T_416,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_418); // @[PositFMA.scala 60:76]
  assign _T_419 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_419); // @[PositFMA.scala 61:33]
  assign _T_420 = sigP[16:0]; // @[PositFMA.scala 62:29]
  assign _T_421 = _T_420 != 17'h0; // @[PositFMA.scala 62:33]
  assign eqTwo = ~ _T_421; // @[PositFMA.scala 62:19]
  assign _T_422 = sigP[18]; // @[PositFMA.scala 64:29]
  assign _T_423 = sigP[17]; // @[PositFMA.scala 64:56]
  assign _T_424 = ~ _T_423; // @[PositFMA.scala 64:51]
  assign _T_425 = _T_422 & _T_424; // @[PositFMA.scala 64:49]
  assign eqFour = _T_425 & eqTwo; // @[PositFMA.scala 64:76]
  assign _T_426 = sigP[19]; // @[PositFMA.scala 66:23]
  assign geTwo = _T_426 ^ _T_423; // @[PositFMA.scala 66:43]
  assign _T_428 = {eqFour,geTwo}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_428)}; // @[PositFMA.scala 67:38]
  assign mulSign = sigP[19:19]; // @[PositFMA.scala 68:28]
  assign _T_429 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 70:30]
  assign _GEN_12 = {{4{expBias[2]}},expBias}; // @[PositFMA.scala 70:44]
  assign _T_431 = $signed(_T_429) + $signed(_GEN_12); // @[PositFMA.scala 70:44]
  assign mulScale = $signed(_T_431); // @[PositFMA.scala 70:44]
  assign _T_432 = sigP[17:0]; // @[PositFMA.scala 73:29]
  assign _T_433 = sigP[16:0]; // @[PositFMA.scala 74:29]
  assign _T_434 = {_T_433, 1'h0}; // @[PositFMA.scala 74:48]
  assign mulSigTmp = geTwo ? _T_432 : _T_434; // @[PositFMA.scala 71:22]
  assign _T_436 = mulSigTmp[17:17]; // @[PositFMA.scala 78:39]
  assign _T_437 = _T_436 | eqFour; // @[PositFMA.scala 78:43]
  assign _T_438 = mulSigTmp[16:0]; // @[PositFMA.scala 79:39]
  assign mulSig = {mulSign,_T_437,_T_438}; // @[Cat.scala 29:58]
  assign _T_464 = ~ addSign_phase2; // @[PositFMA.scala 108:29]
  assign _T_465 = ~ addZero_phase2; // @[PositFMA.scala 108:47]
  assign _T_466 = _T_464 & _T_465; // @[PositFMA.scala 108:45]
  assign extAddSig = {addSign_phase2,_T_466,addFrac_phase2,9'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[5]}},addScale_phase2}; // @[PositFMA.scala 112:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 112:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[5]}},addScale_phase2}); // @[PositFMA.scala 113:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[5]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 114:26]
  assign _T_470 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 115:36]
  assign scaleDiff = $signed(_T_470); // @[PositFMA.scala 115:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 116:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 117:26]
  assign _T_471 = $unsigned(scaleDiff); // @[PositFMA.scala 118:69]
  assign _T_472 = _T_471 < 7'h13; // @[Shift.scala 39:24]
  assign _T_473 = _T_471[4:0]; // @[Shift.scala 40:44]
  assign _T_474 = smallerSigTmp[18:16]; // @[Shift.scala 90:30]
  assign _T_475 = smallerSigTmp[15:0]; // @[Shift.scala 90:48]
  assign _T_476 = _T_475 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{2'd0}, _T_476}; // @[Shift.scala 90:39]
  assign _T_477 = _T_474 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_478 = _T_473[4]; // @[Shift.scala 12:21]
  assign _T_479 = smallerSigTmp[18]; // @[Shift.scala 12:21]
  assign _T_481 = _T_479 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_482 = {_T_481,_T_477}; // @[Cat.scala 29:58]
  assign _T_483 = _T_478 ? _T_482 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_484 = _T_473[3:0]; // @[Shift.scala 92:77]
  assign _T_485 = _T_483[18:8]; // @[Shift.scala 90:30]
  assign _T_486 = _T_483[7:0]; // @[Shift.scala 90:48]
  assign _T_487 = _T_486 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{10'd0}, _T_487}; // @[Shift.scala 90:39]
  assign _T_488 = _T_485 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_489 = _T_484[3]; // @[Shift.scala 12:21]
  assign _T_490 = _T_483[18]; // @[Shift.scala 12:21]
  assign _T_492 = _T_490 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_493 = {_T_492,_T_488}; // @[Cat.scala 29:58]
  assign _T_494 = _T_489 ? _T_493 : _T_483; // @[Shift.scala 91:22]
  assign _T_495 = _T_484[2:0]; // @[Shift.scala 92:77]
  assign _T_496 = _T_494[18:4]; // @[Shift.scala 90:30]
  assign _T_497 = _T_494[3:0]; // @[Shift.scala 90:48]
  assign _T_498 = _T_497 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{14'd0}, _T_498}; // @[Shift.scala 90:39]
  assign _T_499 = _T_496 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_500 = _T_495[2]; // @[Shift.scala 12:21]
  assign _T_501 = _T_494[18]; // @[Shift.scala 12:21]
  assign _T_503 = _T_501 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_504 = {_T_503,_T_499}; // @[Cat.scala 29:58]
  assign _T_505 = _T_500 ? _T_504 : _T_494; // @[Shift.scala 91:22]
  assign _T_506 = _T_495[1:0]; // @[Shift.scala 92:77]
  assign _T_507 = _T_505[18:2]; // @[Shift.scala 90:30]
  assign _T_508 = _T_505[1:0]; // @[Shift.scala 90:48]
  assign _T_509 = _T_508 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_17 = {{16'd0}, _T_509}; // @[Shift.scala 90:39]
  assign _T_510 = _T_507 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_511 = _T_506[1]; // @[Shift.scala 12:21]
  assign _T_512 = _T_505[18]; // @[Shift.scala 12:21]
  assign _T_514 = _T_512 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_515 = {_T_514,_T_510}; // @[Cat.scala 29:58]
  assign _T_516 = _T_511 ? _T_515 : _T_505; // @[Shift.scala 91:22]
  assign _T_517 = _T_506[0:0]; // @[Shift.scala 92:77]
  assign _T_518 = _T_516[18:1]; // @[Shift.scala 90:30]
  assign _T_519 = _T_516[0:0]; // @[Shift.scala 90:48]
  assign _GEN_18 = {{17'd0}, _T_519}; // @[Shift.scala 90:39]
  assign _T_521 = _T_518 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_523 = _T_516[18]; // @[Shift.scala 12:21]
  assign _T_524 = {_T_523,_T_521}; // @[Cat.scala 29:58]
  assign _T_525 = _T_517 ? _T_524 : _T_516; // @[Shift.scala 91:22]
  assign _T_528 = _T_479 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_472 ? _T_525 : _T_528; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 119:34]
  assign _T_529 = mulSig_phase2[18:18]; // @[PositFMA.scala 120:42]
  assign _T_530 = _T_529 ^ addSign_phase2; // @[PositFMA.scala 120:46]
  assign _T_531 = rawSumSig[19:19]; // @[PositFMA.scala 120:79]
  assign sumSign = _T_530 ^ _T_531; // @[PositFMA.scala 120:63]
  assign _T_533 = greaterSig + smallerSig; // @[PositFMA.scala 121:50]
  assign signSumSig = {sumSign,_T_533}; // @[Cat.scala 29:58]
  assign _T_534 = signSumSig[19:1]; // @[PositFMA.scala 125:33]
  assign _T_535 = signSumSig[18:0]; // @[PositFMA.scala 125:68]
  assign sumXor = _T_534 ^ _T_535; // @[PositFMA.scala 125:51]
  assign _T_536 = sumXor[18:3]; // @[LZD.scala 43:32]
  assign _T_537 = _T_536[15:8]; // @[LZD.scala 43:32]
  assign _T_538 = _T_537[7:4]; // @[LZD.scala 43:32]
  assign _T_539 = _T_538[3:2]; // @[LZD.scala 43:32]
  assign _T_540 = _T_539 != 2'h0; // @[LZD.scala 39:14]
  assign _T_541 = _T_539[1]; // @[LZD.scala 39:21]
  assign _T_542 = _T_539[0]; // @[LZD.scala 39:30]
  assign _T_543 = ~ _T_542; // @[LZD.scala 39:27]
  assign _T_544 = _T_541 | _T_543; // @[LZD.scala 39:25]
  assign _T_545 = {_T_540,_T_544}; // @[Cat.scala 29:58]
  assign _T_546 = _T_538[1:0]; // @[LZD.scala 44:32]
  assign _T_547 = _T_546 != 2'h0; // @[LZD.scala 39:14]
  assign _T_548 = _T_546[1]; // @[LZD.scala 39:21]
  assign _T_549 = _T_546[0]; // @[LZD.scala 39:30]
  assign _T_550 = ~ _T_549; // @[LZD.scala 39:27]
  assign _T_551 = _T_548 | _T_550; // @[LZD.scala 39:25]
  assign _T_552 = {_T_547,_T_551}; // @[Cat.scala 29:58]
  assign _T_553 = _T_545[1]; // @[Shift.scala 12:21]
  assign _T_554 = _T_552[1]; // @[Shift.scala 12:21]
  assign _T_555 = _T_553 | _T_554; // @[LZD.scala 49:16]
  assign _T_556 = ~ _T_554; // @[LZD.scala 49:27]
  assign _T_557 = _T_553 | _T_556; // @[LZD.scala 49:25]
  assign _T_558 = _T_545[0:0]; // @[LZD.scala 49:47]
  assign _T_559 = _T_552[0:0]; // @[LZD.scala 49:59]
  assign _T_560 = _T_553 ? _T_558 : _T_559; // @[LZD.scala 49:35]
  assign _T_562 = {_T_555,_T_557,_T_560}; // @[Cat.scala 29:58]
  assign _T_563 = _T_537[3:0]; // @[LZD.scala 44:32]
  assign _T_564 = _T_563[3:2]; // @[LZD.scala 43:32]
  assign _T_565 = _T_564 != 2'h0; // @[LZD.scala 39:14]
  assign _T_566 = _T_564[1]; // @[LZD.scala 39:21]
  assign _T_567 = _T_564[0]; // @[LZD.scala 39:30]
  assign _T_568 = ~ _T_567; // @[LZD.scala 39:27]
  assign _T_569 = _T_566 | _T_568; // @[LZD.scala 39:25]
  assign _T_570 = {_T_565,_T_569}; // @[Cat.scala 29:58]
  assign _T_571 = _T_563[1:0]; // @[LZD.scala 44:32]
  assign _T_572 = _T_571 != 2'h0; // @[LZD.scala 39:14]
  assign _T_573 = _T_571[1]; // @[LZD.scala 39:21]
  assign _T_574 = _T_571[0]; // @[LZD.scala 39:30]
  assign _T_575 = ~ _T_574; // @[LZD.scala 39:27]
  assign _T_576 = _T_573 | _T_575; // @[LZD.scala 39:25]
  assign _T_577 = {_T_572,_T_576}; // @[Cat.scala 29:58]
  assign _T_578 = _T_570[1]; // @[Shift.scala 12:21]
  assign _T_579 = _T_577[1]; // @[Shift.scala 12:21]
  assign _T_580 = _T_578 | _T_579; // @[LZD.scala 49:16]
  assign _T_581 = ~ _T_579; // @[LZD.scala 49:27]
  assign _T_582 = _T_578 | _T_581; // @[LZD.scala 49:25]
  assign _T_583 = _T_570[0:0]; // @[LZD.scala 49:47]
  assign _T_584 = _T_577[0:0]; // @[LZD.scala 49:59]
  assign _T_585 = _T_578 ? _T_583 : _T_584; // @[LZD.scala 49:35]
  assign _T_587 = {_T_580,_T_582,_T_585}; // @[Cat.scala 29:58]
  assign _T_588 = _T_562[2]; // @[Shift.scala 12:21]
  assign _T_589 = _T_587[2]; // @[Shift.scala 12:21]
  assign _T_590 = _T_588 | _T_589; // @[LZD.scala 49:16]
  assign _T_591 = ~ _T_589; // @[LZD.scala 49:27]
  assign _T_592 = _T_588 | _T_591; // @[LZD.scala 49:25]
  assign _T_593 = _T_562[1:0]; // @[LZD.scala 49:47]
  assign _T_594 = _T_587[1:0]; // @[LZD.scala 49:59]
  assign _T_595 = _T_588 ? _T_593 : _T_594; // @[LZD.scala 49:35]
  assign _T_597 = {_T_590,_T_592,_T_595}; // @[Cat.scala 29:58]
  assign _T_598 = _T_536[7:0]; // @[LZD.scala 44:32]
  assign _T_599 = _T_598[7:4]; // @[LZD.scala 43:32]
  assign _T_600 = _T_599[3:2]; // @[LZD.scala 43:32]
  assign _T_601 = _T_600 != 2'h0; // @[LZD.scala 39:14]
  assign _T_602 = _T_600[1]; // @[LZD.scala 39:21]
  assign _T_603 = _T_600[0]; // @[LZD.scala 39:30]
  assign _T_604 = ~ _T_603; // @[LZD.scala 39:27]
  assign _T_605 = _T_602 | _T_604; // @[LZD.scala 39:25]
  assign _T_606 = {_T_601,_T_605}; // @[Cat.scala 29:58]
  assign _T_607 = _T_599[1:0]; // @[LZD.scala 44:32]
  assign _T_608 = _T_607 != 2'h0; // @[LZD.scala 39:14]
  assign _T_609 = _T_607[1]; // @[LZD.scala 39:21]
  assign _T_610 = _T_607[0]; // @[LZD.scala 39:30]
  assign _T_611 = ~ _T_610; // @[LZD.scala 39:27]
  assign _T_612 = _T_609 | _T_611; // @[LZD.scala 39:25]
  assign _T_613 = {_T_608,_T_612}; // @[Cat.scala 29:58]
  assign _T_614 = _T_606[1]; // @[Shift.scala 12:21]
  assign _T_615 = _T_613[1]; // @[Shift.scala 12:21]
  assign _T_616 = _T_614 | _T_615; // @[LZD.scala 49:16]
  assign _T_617 = ~ _T_615; // @[LZD.scala 49:27]
  assign _T_618 = _T_614 | _T_617; // @[LZD.scala 49:25]
  assign _T_619 = _T_606[0:0]; // @[LZD.scala 49:47]
  assign _T_620 = _T_613[0:0]; // @[LZD.scala 49:59]
  assign _T_621 = _T_614 ? _T_619 : _T_620; // @[LZD.scala 49:35]
  assign _T_623 = {_T_616,_T_618,_T_621}; // @[Cat.scala 29:58]
  assign _T_624 = _T_598[3:0]; // @[LZD.scala 44:32]
  assign _T_625 = _T_624[3:2]; // @[LZD.scala 43:32]
  assign _T_626 = _T_625 != 2'h0; // @[LZD.scala 39:14]
  assign _T_627 = _T_625[1]; // @[LZD.scala 39:21]
  assign _T_628 = _T_625[0]; // @[LZD.scala 39:30]
  assign _T_629 = ~ _T_628; // @[LZD.scala 39:27]
  assign _T_630 = _T_627 | _T_629; // @[LZD.scala 39:25]
  assign _T_631 = {_T_626,_T_630}; // @[Cat.scala 29:58]
  assign _T_632 = _T_624[1:0]; // @[LZD.scala 44:32]
  assign _T_633 = _T_632 != 2'h0; // @[LZD.scala 39:14]
  assign _T_634 = _T_632[1]; // @[LZD.scala 39:21]
  assign _T_635 = _T_632[0]; // @[LZD.scala 39:30]
  assign _T_636 = ~ _T_635; // @[LZD.scala 39:27]
  assign _T_637 = _T_634 | _T_636; // @[LZD.scala 39:25]
  assign _T_638 = {_T_633,_T_637}; // @[Cat.scala 29:58]
  assign _T_639 = _T_631[1]; // @[Shift.scala 12:21]
  assign _T_640 = _T_638[1]; // @[Shift.scala 12:21]
  assign _T_641 = _T_639 | _T_640; // @[LZD.scala 49:16]
  assign _T_642 = ~ _T_640; // @[LZD.scala 49:27]
  assign _T_643 = _T_639 | _T_642; // @[LZD.scala 49:25]
  assign _T_644 = _T_631[0:0]; // @[LZD.scala 49:47]
  assign _T_645 = _T_638[0:0]; // @[LZD.scala 49:59]
  assign _T_646 = _T_639 ? _T_644 : _T_645; // @[LZD.scala 49:35]
  assign _T_648 = {_T_641,_T_643,_T_646}; // @[Cat.scala 29:58]
  assign _T_649 = _T_623[2]; // @[Shift.scala 12:21]
  assign _T_650 = _T_648[2]; // @[Shift.scala 12:21]
  assign _T_651 = _T_649 | _T_650; // @[LZD.scala 49:16]
  assign _T_652 = ~ _T_650; // @[LZD.scala 49:27]
  assign _T_653 = _T_649 | _T_652; // @[LZD.scala 49:25]
  assign _T_654 = _T_623[1:0]; // @[LZD.scala 49:47]
  assign _T_655 = _T_648[1:0]; // @[LZD.scala 49:59]
  assign _T_656 = _T_649 ? _T_654 : _T_655; // @[LZD.scala 49:35]
  assign _T_658 = {_T_651,_T_653,_T_656}; // @[Cat.scala 29:58]
  assign _T_659 = _T_597[3]; // @[Shift.scala 12:21]
  assign _T_660 = _T_658[3]; // @[Shift.scala 12:21]
  assign _T_661 = _T_659 | _T_660; // @[LZD.scala 49:16]
  assign _T_662 = ~ _T_660; // @[LZD.scala 49:27]
  assign _T_663 = _T_659 | _T_662; // @[LZD.scala 49:25]
  assign _T_664 = _T_597[2:0]; // @[LZD.scala 49:47]
  assign _T_665 = _T_658[2:0]; // @[LZD.scala 49:59]
  assign _T_666 = _T_659 ? _T_664 : _T_665; // @[LZD.scala 49:35]
  assign _T_668 = {_T_661,_T_663,_T_666}; // @[Cat.scala 29:58]
  assign _T_669 = sumXor[2:0]; // @[LZD.scala 44:32]
  assign _T_670 = _T_669[2:1]; // @[LZD.scala 43:32]
  assign _T_671 = _T_670 != 2'h0; // @[LZD.scala 39:14]
  assign _T_672 = _T_670[1]; // @[LZD.scala 39:21]
  assign _T_673 = _T_670[0]; // @[LZD.scala 39:30]
  assign _T_674 = ~ _T_673; // @[LZD.scala 39:27]
  assign _T_675 = _T_672 | _T_674; // @[LZD.scala 39:25]
  assign _T_676 = {_T_671,_T_675}; // @[Cat.scala 29:58]
  assign _T_677 = _T_669[0:0]; // @[LZD.scala 44:32]
  assign _T_679 = _T_676[1]; // @[Shift.scala 12:21]
  assign _T_681 = _T_676[0:0]; // @[LZD.scala 55:32]
  assign _T_682 = _T_679 ? _T_681 : _T_677; // @[LZD.scala 55:20]
  assign _T_684 = _T_668[4]; // @[Shift.scala 12:21]
  assign _T_687 = {2'h3,_T_679,_T_682}; // @[Cat.scala 29:58]
  assign _T_688 = _T_668[3:0]; // @[LZD.scala 55:32]
  assign _T_689 = _T_684 ? _T_688 : _T_687; // @[LZD.scala 55:20]
  assign sumLZD = {_T_684,_T_689}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 127:24]
  assign _T_690 = signSumSig[17:0]; // @[PositFMA.scala 128:38]
  assign _T_691 = shiftValue < 5'h12; // @[Shift.scala 16:24]
  assign _T_693 = shiftValue[4]; // @[Shift.scala 12:21]
  assign _T_694 = _T_690[1:0]; // @[Shift.scala 64:52]
  assign _T_696 = {_T_694,16'h0}; // @[Cat.scala 29:58]
  assign _T_697 = _T_693 ? _T_696 : _T_690; // @[Shift.scala 64:27]
  assign _T_698 = shiftValue[3:0]; // @[Shift.scala 66:70]
  assign _T_699 = _T_698[3]; // @[Shift.scala 12:21]
  assign _T_700 = _T_697[9:0]; // @[Shift.scala 64:52]
  assign _T_702 = {_T_700,8'h0}; // @[Cat.scala 29:58]
  assign _T_703 = _T_699 ? _T_702 : _T_697; // @[Shift.scala 64:27]
  assign _T_704 = _T_698[2:0]; // @[Shift.scala 66:70]
  assign _T_705 = _T_704[2]; // @[Shift.scala 12:21]
  assign _T_706 = _T_703[13:0]; // @[Shift.scala 64:52]
  assign _T_708 = {_T_706,4'h0}; // @[Cat.scala 29:58]
  assign _T_709 = _T_705 ? _T_708 : _T_703; // @[Shift.scala 64:27]
  assign _T_710 = _T_704[1:0]; // @[Shift.scala 66:70]
  assign _T_711 = _T_710[1]; // @[Shift.scala 12:21]
  assign _T_712 = _T_709[15:0]; // @[Shift.scala 64:52]
  assign _T_714 = {_T_712,2'h0}; // @[Cat.scala 29:58]
  assign _T_715 = _T_711 ? _T_714 : _T_709; // @[Shift.scala 64:27]
  assign _T_716 = _T_710[0:0]; // @[Shift.scala 66:70]
  assign _T_718 = _T_715[16:0]; // @[Shift.scala 64:52]
  assign _T_719 = {_T_718,1'h0}; // @[Cat.scala 29:58]
  assign _T_720 = _T_716 ? _T_719 : _T_715; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_691 ? _T_720 : 18'h0; // @[Shift.scala 16:10]
  assign _T_722 = $signed(greaterScale) + $signed(7'sh2); // @[PositFMA.scala 131:36]
  assign _T_723 = $signed(_T_722); // @[PositFMA.scala 131:36]
  assign _T_724 = {1'h1,_T_684,_T_689}; // @[Cat.scala 29:58]
  assign _T_725 = $signed(_T_724); // @[PositFMA.scala 131:61]
  assign _GEN_19 = {{1{_T_725[5]}},_T_725}; // @[PositFMA.scala 131:42]
  assign _T_727 = $signed(_T_723) + $signed(_GEN_19); // @[PositFMA.scala 131:42]
  assign sumScale = $signed(_T_727); // @[PositFMA.scala 131:42]
  assign sumFrac = normalFracTmp[17:10]; // @[PositFMA.scala 132:41]
  assign grsTmp = normalFracTmp[9:0]; // @[PositFMA.scala 135:41]
  assign _T_728 = grsTmp[9:8]; // @[PositFMA.scala 138:40]
  assign _T_729 = grsTmp[7:0]; // @[PositFMA.scala 138:56]
  assign _T_730 = _T_729 != 8'h0; // @[PositFMA.scala 138:60]
  assign underflow = $signed(sumScale) < $signed(-7'sh14); // @[PositFMA.scala 145:32]
  assign overflow = $signed(sumScale) > $signed(7'sh14); // @[PositFMA.scala 146:32]
  assign _T_731 = signSumSig != 20'h0; // @[PositFMA.scala 155:32]
  assign decF_isZero = ~ _T_731; // @[PositFMA.scala 155:20]
  assign _T_733 = underflow ? $signed(-7'sh14) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_734 = overflow ? $signed(7'sh14) : $signed(_T_733); // @[Mux.scala 87:16]
  assign _GEN_20 = _T_734[5:0]; // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  assign decF_scale = $signed(_GEN_20); // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  assign _T_735 = decF_scale[0]; // @[convert.scala 46:61]
  assign _T_736 = ~ _T_735; // @[convert.scala 46:52]
  assign _T_738 = sumSign ? _T_736 : _T_735; // @[convert.scala 46:42]
  assign _T_739 = decF_scale[5:1]; // @[convert.scala 48:34]
  assign _T_740 = _T_739[4:4]; // @[convert.scala 49:36]
  assign _T_742 = ~ _T_739; // @[convert.scala 50:36]
  assign _T_743 = $signed(_T_742); // @[convert.scala 50:36]
  assign _T_744 = _T_740 ? $signed(_T_743) : $signed(_T_739); // @[convert.scala 50:28]
  assign _T_745 = _T_740 ^ sumSign; // @[convert.scala 51:31]
  assign _T_746 = ~ _T_745; // @[convert.scala 52:43]
  assign _T_750 = {_T_746,_T_745,_T_738,sumFrac,_T_728,_T_730}; // @[Cat.scala 29:58]
  assign _T_751 = $unsigned(_T_744); // @[Shift.scala 39:17]
  assign _T_752 = _T_751 < 5'he; // @[Shift.scala 39:24]
  assign _T_753 = _T_744[3:0]; // @[Shift.scala 40:44]
  assign _T_754 = _T_750[13:8]; // @[Shift.scala 90:30]
  assign _T_755 = _T_750[7:0]; // @[Shift.scala 90:48]
  assign _T_756 = _T_755 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{5'd0}, _T_756}; // @[Shift.scala 90:39]
  assign _T_757 = _T_754 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_758 = _T_753[3]; // @[Shift.scala 12:21]
  assign _T_759 = _T_750[13]; // @[Shift.scala 12:21]
  assign _T_761 = _T_759 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_762 = {_T_761,_T_757}; // @[Cat.scala 29:58]
  assign _T_763 = _T_758 ? _T_762 : _T_750; // @[Shift.scala 91:22]
  assign _T_764 = _T_753[2:0]; // @[Shift.scala 92:77]
  assign _T_765 = _T_763[13:4]; // @[Shift.scala 90:30]
  assign _T_766 = _T_763[3:0]; // @[Shift.scala 90:48]
  assign _T_767 = _T_766 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{9'd0}, _T_767}; // @[Shift.scala 90:39]
  assign _T_768 = _T_765 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_769 = _T_764[2]; // @[Shift.scala 12:21]
  assign _T_770 = _T_763[13]; // @[Shift.scala 12:21]
  assign _T_772 = _T_770 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_773 = {_T_772,_T_768}; // @[Cat.scala 29:58]
  assign _T_774 = _T_769 ? _T_773 : _T_763; // @[Shift.scala 91:22]
  assign _T_775 = _T_764[1:0]; // @[Shift.scala 92:77]
  assign _T_776 = _T_774[13:2]; // @[Shift.scala 90:30]
  assign _T_777 = _T_774[1:0]; // @[Shift.scala 90:48]
  assign _T_778 = _T_777 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{11'd0}, _T_778}; // @[Shift.scala 90:39]
  assign _T_779 = _T_776 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_780 = _T_775[1]; // @[Shift.scala 12:21]
  assign _T_781 = _T_774[13]; // @[Shift.scala 12:21]
  assign _T_783 = _T_781 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_784 = {_T_783,_T_779}; // @[Cat.scala 29:58]
  assign _T_785 = _T_780 ? _T_784 : _T_774; // @[Shift.scala 91:22]
  assign _T_786 = _T_775[0:0]; // @[Shift.scala 92:77]
  assign _T_787 = _T_785[13:1]; // @[Shift.scala 90:30]
  assign _T_788 = _T_785[0:0]; // @[Shift.scala 90:48]
  assign _GEN_24 = {{12'd0}, _T_788}; // @[Shift.scala 90:39]
  assign _T_790 = _T_787 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_792 = _T_785[13]; // @[Shift.scala 12:21]
  assign _T_793 = {_T_792,_T_790}; // @[Cat.scala 29:58]
  assign _T_794 = _T_786 ? _T_793 : _T_785; // @[Shift.scala 91:22]
  assign _T_797 = _T_759 ? 14'h3fff : 14'h0; // @[Bitwise.scala 71:12]
  assign _T_798 = _T_752 ? _T_794 : _T_797; // @[Shift.scala 39:10]
  assign _T_799 = _T_798[3]; // @[convert.scala 55:31]
  assign _T_800 = _T_798[2]; // @[convert.scala 56:31]
  assign _T_801 = _T_798[1]; // @[convert.scala 57:31]
  assign _T_802 = _T_798[0]; // @[convert.scala 58:31]
  assign _T_803 = _T_798[13:3]; // @[convert.scala 59:69]
  assign _T_804 = _T_803 != 11'h0; // @[convert.scala 59:81]
  assign _T_805 = ~ _T_804; // @[convert.scala 59:50]
  assign _T_807 = _T_803 == 11'h7ff; // @[convert.scala 60:81]
  assign _T_808 = _T_799 | _T_801; // @[convert.scala 61:44]
  assign _T_809 = _T_808 | _T_802; // @[convert.scala 61:52]
  assign _T_810 = _T_800 & _T_809; // @[convert.scala 61:36]
  assign _T_811 = ~ _T_807; // @[convert.scala 62:63]
  assign _T_812 = _T_811 & _T_810; // @[convert.scala 62:103]
  assign _T_813 = _T_805 | _T_812; // @[convert.scala 62:60]
  assign _GEN_25 = {{10'd0}, _T_813}; // @[convert.scala 63:56]
  assign _T_816 = _T_803 + _GEN_25; // @[convert.scala 63:56]
  assign _T_817 = {sumSign,_T_816}; // @[Cat.scala 29:58]
  assign io_F = _T_825; // @[PositFMA.scala 175:15]
  assign io_outValid = _T_821; // @[PositFMA.scala 174:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_821 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_825 = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_277;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_821 <= 1'h0;
    end else begin
      _T_821 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_825 <= 12'h800;
      end else begin
        if (decF_isZero) begin
          _T_825 <= 12'h0;
        end else begin
          _T_825 <= _T_817;
        end
      end
    end
  end
endmodule
