module PositFMA29_3(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [1:0]  io_fmaOp,
  input  [28:0] io_A,
  input  [28:0] io_B,
  input  [28:0] io_C,
  output [28:0] io_F,
  output        io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [28:0] _T_2; // @[Bitwise.scala 71:12]
  wire [28:0] _T_3; // @[PositFMA.scala 47:41]
  wire [28:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [28:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [28:0] _T_8; // @[Bitwise.scala 71:12]
  wire [28:0] _T_9; // @[PositFMA.scala 48:41]
  wire [28:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [28:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [26:0] _T_16; // @[convert.scala 19:24]
  wire [26:0] _T_17; // @[convert.scala 19:43]
  wire [26:0] _T_18; // @[convert.scala 19:39]
  wire [15:0] _T_19; // @[LZD.scala 43:32]
  wire [7:0] _T_20; // @[LZD.scala 43:32]
  wire [3:0] _T_21; // @[LZD.scala 43:32]
  wire [1:0] _T_22; // @[LZD.scala 43:32]
  wire  _T_23; // @[LZD.scala 39:14]
  wire  _T_24; // @[LZD.scala 39:21]
  wire  _T_25; // @[LZD.scala 39:30]
  wire  _T_26; // @[LZD.scala 39:27]
  wire  _T_27; // @[LZD.scala 39:25]
  wire [1:0] _T_28; // @[Cat.scala 29:58]
  wire [1:0] _T_29; // @[LZD.scala 44:32]
  wire  _T_30; // @[LZD.scala 39:14]
  wire  _T_31; // @[LZD.scala 39:21]
  wire  _T_32; // @[LZD.scala 39:30]
  wire  _T_33; // @[LZD.scala 39:27]
  wire  _T_34; // @[LZD.scala 39:25]
  wire [1:0] _T_35; // @[Cat.scala 29:58]
  wire  _T_36; // @[Shift.scala 12:21]
  wire  _T_37; // @[Shift.scala 12:21]
  wire  _T_38; // @[LZD.scala 49:16]
  wire  _T_39; // @[LZD.scala 49:27]
  wire  _T_40; // @[LZD.scala 49:25]
  wire  _T_41; // @[LZD.scala 49:47]
  wire  _T_42; // @[LZD.scala 49:59]
  wire  _T_43; // @[LZD.scala 49:35]
  wire [2:0] _T_45; // @[Cat.scala 29:58]
  wire [3:0] _T_46; // @[LZD.scala 44:32]
  wire [1:0] _T_47; // @[LZD.scala 43:32]
  wire  _T_48; // @[LZD.scala 39:14]
  wire  _T_49; // @[LZD.scala 39:21]
  wire  _T_50; // @[LZD.scala 39:30]
  wire  _T_51; // @[LZD.scala 39:27]
  wire  _T_52; // @[LZD.scala 39:25]
  wire [1:0] _T_53; // @[Cat.scala 29:58]
  wire [1:0] _T_54; // @[LZD.scala 44:32]
  wire  _T_55; // @[LZD.scala 39:14]
  wire  _T_56; // @[LZD.scala 39:21]
  wire  _T_57; // @[LZD.scala 39:30]
  wire  _T_58; // @[LZD.scala 39:27]
  wire  _T_59; // @[LZD.scala 39:25]
  wire [1:0] _T_60; // @[Cat.scala 29:58]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[Shift.scala 12:21]
  wire  _T_63; // @[LZD.scala 49:16]
  wire  _T_64; // @[LZD.scala 49:27]
  wire  _T_65; // @[LZD.scala 49:25]
  wire  _T_66; // @[LZD.scala 49:47]
  wire  _T_67; // @[LZD.scala 49:59]
  wire  _T_68; // @[LZD.scala 49:35]
  wire [2:0] _T_70; // @[Cat.scala 29:58]
  wire  _T_71; // @[Shift.scala 12:21]
  wire  _T_72; // @[Shift.scala 12:21]
  wire  _T_73; // @[LZD.scala 49:16]
  wire  _T_74; // @[LZD.scala 49:27]
  wire  _T_75; // @[LZD.scala 49:25]
  wire [1:0] _T_76; // @[LZD.scala 49:47]
  wire [1:0] _T_77; // @[LZD.scala 49:59]
  wire [1:0] _T_78; // @[LZD.scala 49:35]
  wire [3:0] _T_80; // @[Cat.scala 29:58]
  wire [7:0] _T_81; // @[LZD.scala 44:32]
  wire [3:0] _T_82; // @[LZD.scala 43:32]
  wire [1:0] _T_83; // @[LZD.scala 43:32]
  wire  _T_84; // @[LZD.scala 39:14]
  wire  _T_85; // @[LZD.scala 39:21]
  wire  _T_86; // @[LZD.scala 39:30]
  wire  _T_87; // @[LZD.scala 39:27]
  wire  _T_88; // @[LZD.scala 39:25]
  wire [1:0] _T_89; // @[Cat.scala 29:58]
  wire [1:0] _T_90; // @[LZD.scala 44:32]
  wire  _T_91; // @[LZD.scala 39:14]
  wire  _T_92; // @[LZD.scala 39:21]
  wire  _T_93; // @[LZD.scala 39:30]
  wire  _T_94; // @[LZD.scala 39:27]
  wire  _T_95; // @[LZD.scala 39:25]
  wire [1:0] _T_96; // @[Cat.scala 29:58]
  wire  _T_97; // @[Shift.scala 12:21]
  wire  _T_98; // @[Shift.scala 12:21]
  wire  _T_99; // @[LZD.scala 49:16]
  wire  _T_100; // @[LZD.scala 49:27]
  wire  _T_101; // @[LZD.scala 49:25]
  wire  _T_102; // @[LZD.scala 49:47]
  wire  _T_103; // @[LZD.scala 49:59]
  wire  _T_104; // @[LZD.scala 49:35]
  wire [2:0] _T_106; // @[Cat.scala 29:58]
  wire [3:0] _T_107; // @[LZD.scala 44:32]
  wire [1:0] _T_108; // @[LZD.scala 43:32]
  wire  _T_109; // @[LZD.scala 39:14]
  wire  _T_110; // @[LZD.scala 39:21]
  wire  _T_111; // @[LZD.scala 39:30]
  wire  _T_112; // @[LZD.scala 39:27]
  wire  _T_113; // @[LZD.scala 39:25]
  wire [1:0] _T_114; // @[Cat.scala 29:58]
  wire [1:0] _T_115; // @[LZD.scala 44:32]
  wire  _T_116; // @[LZD.scala 39:14]
  wire  _T_117; // @[LZD.scala 39:21]
  wire  _T_118; // @[LZD.scala 39:30]
  wire  _T_119; // @[LZD.scala 39:27]
  wire  _T_120; // @[LZD.scala 39:25]
  wire [1:0] _T_121; // @[Cat.scala 29:58]
  wire  _T_122; // @[Shift.scala 12:21]
  wire  _T_123; // @[Shift.scala 12:21]
  wire  _T_124; // @[LZD.scala 49:16]
  wire  _T_125; // @[LZD.scala 49:27]
  wire  _T_126; // @[LZD.scala 49:25]
  wire  _T_127; // @[LZD.scala 49:47]
  wire  _T_128; // @[LZD.scala 49:59]
  wire  _T_129; // @[LZD.scala 49:35]
  wire [2:0] _T_131; // @[Cat.scala 29:58]
  wire  _T_132; // @[Shift.scala 12:21]
  wire  _T_133; // @[Shift.scala 12:21]
  wire  _T_134; // @[LZD.scala 49:16]
  wire  _T_135; // @[LZD.scala 49:27]
  wire  _T_136; // @[LZD.scala 49:25]
  wire [1:0] _T_137; // @[LZD.scala 49:47]
  wire [1:0] _T_138; // @[LZD.scala 49:59]
  wire [1:0] _T_139; // @[LZD.scala 49:35]
  wire [3:0] _T_141; // @[Cat.scala 29:58]
  wire  _T_142; // @[Shift.scala 12:21]
  wire  _T_143; // @[Shift.scala 12:21]
  wire  _T_144; // @[LZD.scala 49:16]
  wire  _T_145; // @[LZD.scala 49:27]
  wire  _T_146; // @[LZD.scala 49:25]
  wire [2:0] _T_147; // @[LZD.scala 49:47]
  wire [2:0] _T_148; // @[LZD.scala 49:59]
  wire [2:0] _T_149; // @[LZD.scala 49:35]
  wire [4:0] _T_151; // @[Cat.scala 29:58]
  wire [10:0] _T_152; // @[LZD.scala 44:32]
  wire [7:0] _T_153; // @[LZD.scala 43:32]
  wire [3:0] _T_154; // @[LZD.scala 43:32]
  wire [1:0] _T_155; // @[LZD.scala 43:32]
  wire  _T_156; // @[LZD.scala 39:14]
  wire  _T_157; // @[LZD.scala 39:21]
  wire  _T_158; // @[LZD.scala 39:30]
  wire  _T_159; // @[LZD.scala 39:27]
  wire  _T_160; // @[LZD.scala 39:25]
  wire [1:0] _T_161; // @[Cat.scala 29:58]
  wire [1:0] _T_162; // @[LZD.scala 44:32]
  wire  _T_163; // @[LZD.scala 39:14]
  wire  _T_164; // @[LZD.scala 39:21]
  wire  _T_165; // @[LZD.scala 39:30]
  wire  _T_166; // @[LZD.scala 39:27]
  wire  _T_167; // @[LZD.scala 39:25]
  wire [1:0] _T_168; // @[Cat.scala 29:58]
  wire  _T_169; // @[Shift.scala 12:21]
  wire  _T_170; // @[Shift.scala 12:21]
  wire  _T_171; // @[LZD.scala 49:16]
  wire  _T_172; // @[LZD.scala 49:27]
  wire  _T_173; // @[LZD.scala 49:25]
  wire  _T_174; // @[LZD.scala 49:47]
  wire  _T_175; // @[LZD.scala 49:59]
  wire  _T_176; // @[LZD.scala 49:35]
  wire [2:0] _T_178; // @[Cat.scala 29:58]
  wire [3:0] _T_179; // @[LZD.scala 44:32]
  wire [1:0] _T_180; // @[LZD.scala 43:32]
  wire  _T_181; // @[LZD.scala 39:14]
  wire  _T_182; // @[LZD.scala 39:21]
  wire  _T_183; // @[LZD.scala 39:30]
  wire  _T_184; // @[LZD.scala 39:27]
  wire  _T_185; // @[LZD.scala 39:25]
  wire [1:0] _T_186; // @[Cat.scala 29:58]
  wire [1:0] _T_187; // @[LZD.scala 44:32]
  wire  _T_188; // @[LZD.scala 39:14]
  wire  _T_189; // @[LZD.scala 39:21]
  wire  _T_190; // @[LZD.scala 39:30]
  wire  _T_191; // @[LZD.scala 39:27]
  wire  _T_192; // @[LZD.scala 39:25]
  wire [1:0] _T_193; // @[Cat.scala 29:58]
  wire  _T_194; // @[Shift.scala 12:21]
  wire  _T_195; // @[Shift.scala 12:21]
  wire  _T_196; // @[LZD.scala 49:16]
  wire  _T_197; // @[LZD.scala 49:27]
  wire  _T_198; // @[LZD.scala 49:25]
  wire  _T_199; // @[LZD.scala 49:47]
  wire  _T_200; // @[LZD.scala 49:59]
  wire  _T_201; // @[LZD.scala 49:35]
  wire [2:0] _T_203; // @[Cat.scala 29:58]
  wire  _T_204; // @[Shift.scala 12:21]
  wire  _T_205; // @[Shift.scala 12:21]
  wire  _T_206; // @[LZD.scala 49:16]
  wire  _T_207; // @[LZD.scala 49:27]
  wire  _T_208; // @[LZD.scala 49:25]
  wire [1:0] _T_209; // @[LZD.scala 49:47]
  wire [1:0] _T_210; // @[LZD.scala 49:59]
  wire [1:0] _T_211; // @[LZD.scala 49:35]
  wire [3:0] _T_213; // @[Cat.scala 29:58]
  wire [2:0] _T_214; // @[LZD.scala 44:32]
  wire [1:0] _T_215; // @[LZD.scala 43:32]
  wire  _T_216; // @[LZD.scala 39:14]
  wire  _T_217; // @[LZD.scala 39:21]
  wire  _T_218; // @[LZD.scala 39:30]
  wire  _T_219; // @[LZD.scala 39:27]
  wire  _T_220; // @[LZD.scala 39:25]
  wire [1:0] _T_221; // @[Cat.scala 29:58]
  wire  _T_222; // @[LZD.scala 44:32]
  wire  _T_224; // @[Shift.scala 12:21]
  wire  _T_226; // @[LZD.scala 55:32]
  wire  _T_227; // @[LZD.scala 55:20]
  wire  _T_229; // @[Shift.scala 12:21]
  wire [2:0] _T_231; // @[Cat.scala 29:58]
  wire [2:0] _T_232; // @[LZD.scala 55:32]
  wire [2:0] _T_233; // @[LZD.scala 55:20]
  wire [3:0] _T_234; // @[Cat.scala 29:58]
  wire  _T_235; // @[Shift.scala 12:21]
  wire [3:0] _T_237; // @[LZD.scala 55:32]
  wire [3:0] _T_238; // @[LZD.scala 55:20]
  wire [4:0] _T_239; // @[Cat.scala 29:58]
  wire [4:0] _T_240; // @[convert.scala 21:22]
  wire [25:0] _T_241; // @[convert.scala 22:36]
  wire  _T_242; // @[Shift.scala 16:24]
  wire  _T_244; // @[Shift.scala 12:21]
  wire [9:0] _T_245; // @[Shift.scala 64:52]
  wire [25:0] _T_247; // @[Cat.scala 29:58]
  wire [25:0] _T_248; // @[Shift.scala 64:27]
  wire [3:0] _T_249; // @[Shift.scala 66:70]
  wire  _T_250; // @[Shift.scala 12:21]
  wire [17:0] _T_251; // @[Shift.scala 64:52]
  wire [25:0] _T_253; // @[Cat.scala 29:58]
  wire [25:0] _T_254; // @[Shift.scala 64:27]
  wire [2:0] _T_255; // @[Shift.scala 66:70]
  wire  _T_256; // @[Shift.scala 12:21]
  wire [21:0] _T_257; // @[Shift.scala 64:52]
  wire [25:0] _T_259; // @[Cat.scala 29:58]
  wire [25:0] _T_260; // @[Shift.scala 64:27]
  wire [1:0] _T_261; // @[Shift.scala 66:70]
  wire  _T_262; // @[Shift.scala 12:21]
  wire [23:0] _T_263; // @[Shift.scala 64:52]
  wire [25:0] _T_265; // @[Cat.scala 29:58]
  wire [25:0] _T_266; // @[Shift.scala 64:27]
  wire  _T_267; // @[Shift.scala 66:70]
  wire [24:0] _T_269; // @[Shift.scala 64:52]
  wire [25:0] _T_270; // @[Cat.scala 29:58]
  wire [25:0] _T_271; // @[Shift.scala 64:27]
  wire [25:0] _T_272; // @[Shift.scala 16:10]
  wire [2:0] _T_273; // @[convert.scala 23:34]
  wire [22:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_275; // @[convert.scala 25:26]
  wire [4:0] _T_277; // @[convert.scala 25:42]
  wire [2:0] _T_280; // @[convert.scala 26:67]
  wire [2:0] _T_281; // @[convert.scala 26:51]
  wire [8:0] _T_282; // @[Cat.scala 29:58]
  wire [27:0] _T_284; // @[convert.scala 29:56]
  wire  _T_285; // @[convert.scala 29:60]
  wire  _T_286; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_289; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [8:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_298; // @[convert.scala 18:24]
  wire  _T_299; // @[convert.scala 18:40]
  wire  _T_300; // @[convert.scala 18:36]
  wire [26:0] _T_301; // @[convert.scala 19:24]
  wire [26:0] _T_302; // @[convert.scala 19:43]
  wire [26:0] _T_303; // @[convert.scala 19:39]
  wire [15:0] _T_304; // @[LZD.scala 43:32]
  wire [7:0] _T_305; // @[LZD.scala 43:32]
  wire [3:0] _T_306; // @[LZD.scala 43:32]
  wire [1:0] _T_307; // @[LZD.scala 43:32]
  wire  _T_308; // @[LZD.scala 39:14]
  wire  _T_309; // @[LZD.scala 39:21]
  wire  _T_310; // @[LZD.scala 39:30]
  wire  _T_311; // @[LZD.scala 39:27]
  wire  _T_312; // @[LZD.scala 39:25]
  wire [1:0] _T_313; // @[Cat.scala 29:58]
  wire [1:0] _T_314; // @[LZD.scala 44:32]
  wire  _T_315; // @[LZD.scala 39:14]
  wire  _T_316; // @[LZD.scala 39:21]
  wire  _T_317; // @[LZD.scala 39:30]
  wire  _T_318; // @[LZD.scala 39:27]
  wire  _T_319; // @[LZD.scala 39:25]
  wire [1:0] _T_320; // @[Cat.scala 29:58]
  wire  _T_321; // @[Shift.scala 12:21]
  wire  _T_322; // @[Shift.scala 12:21]
  wire  _T_323; // @[LZD.scala 49:16]
  wire  _T_324; // @[LZD.scala 49:27]
  wire  _T_325; // @[LZD.scala 49:25]
  wire  _T_326; // @[LZD.scala 49:47]
  wire  _T_327; // @[LZD.scala 49:59]
  wire  _T_328; // @[LZD.scala 49:35]
  wire [2:0] _T_330; // @[Cat.scala 29:58]
  wire [3:0] _T_331; // @[LZD.scala 44:32]
  wire [1:0] _T_332; // @[LZD.scala 43:32]
  wire  _T_333; // @[LZD.scala 39:14]
  wire  _T_334; // @[LZD.scala 39:21]
  wire  _T_335; // @[LZD.scala 39:30]
  wire  _T_336; // @[LZD.scala 39:27]
  wire  _T_337; // @[LZD.scala 39:25]
  wire [1:0] _T_338; // @[Cat.scala 29:58]
  wire [1:0] _T_339; // @[LZD.scala 44:32]
  wire  _T_340; // @[LZD.scala 39:14]
  wire  _T_341; // @[LZD.scala 39:21]
  wire  _T_342; // @[LZD.scala 39:30]
  wire  _T_343; // @[LZD.scala 39:27]
  wire  _T_344; // @[LZD.scala 39:25]
  wire [1:0] _T_345; // @[Cat.scala 29:58]
  wire  _T_346; // @[Shift.scala 12:21]
  wire  _T_347; // @[Shift.scala 12:21]
  wire  _T_348; // @[LZD.scala 49:16]
  wire  _T_349; // @[LZD.scala 49:27]
  wire  _T_350; // @[LZD.scala 49:25]
  wire  _T_351; // @[LZD.scala 49:47]
  wire  _T_352; // @[LZD.scala 49:59]
  wire  _T_353; // @[LZD.scala 49:35]
  wire [2:0] _T_355; // @[Cat.scala 29:58]
  wire  _T_356; // @[Shift.scala 12:21]
  wire  _T_357; // @[Shift.scala 12:21]
  wire  _T_358; // @[LZD.scala 49:16]
  wire  _T_359; // @[LZD.scala 49:27]
  wire  _T_360; // @[LZD.scala 49:25]
  wire [1:0] _T_361; // @[LZD.scala 49:47]
  wire [1:0] _T_362; // @[LZD.scala 49:59]
  wire [1:0] _T_363; // @[LZD.scala 49:35]
  wire [3:0] _T_365; // @[Cat.scala 29:58]
  wire [7:0] _T_366; // @[LZD.scala 44:32]
  wire [3:0] _T_367; // @[LZD.scala 43:32]
  wire [1:0] _T_368; // @[LZD.scala 43:32]
  wire  _T_369; // @[LZD.scala 39:14]
  wire  _T_370; // @[LZD.scala 39:21]
  wire  _T_371; // @[LZD.scala 39:30]
  wire  _T_372; // @[LZD.scala 39:27]
  wire  _T_373; // @[LZD.scala 39:25]
  wire [1:0] _T_374; // @[Cat.scala 29:58]
  wire [1:0] _T_375; // @[LZD.scala 44:32]
  wire  _T_376; // @[LZD.scala 39:14]
  wire  _T_377; // @[LZD.scala 39:21]
  wire  _T_378; // @[LZD.scala 39:30]
  wire  _T_379; // @[LZD.scala 39:27]
  wire  _T_380; // @[LZD.scala 39:25]
  wire [1:0] _T_381; // @[Cat.scala 29:58]
  wire  _T_382; // @[Shift.scala 12:21]
  wire  _T_383; // @[Shift.scala 12:21]
  wire  _T_384; // @[LZD.scala 49:16]
  wire  _T_385; // @[LZD.scala 49:27]
  wire  _T_386; // @[LZD.scala 49:25]
  wire  _T_387; // @[LZD.scala 49:47]
  wire  _T_388; // @[LZD.scala 49:59]
  wire  _T_389; // @[LZD.scala 49:35]
  wire [2:0] _T_391; // @[Cat.scala 29:58]
  wire [3:0] _T_392; // @[LZD.scala 44:32]
  wire [1:0] _T_393; // @[LZD.scala 43:32]
  wire  _T_394; // @[LZD.scala 39:14]
  wire  _T_395; // @[LZD.scala 39:21]
  wire  _T_396; // @[LZD.scala 39:30]
  wire  _T_397; // @[LZD.scala 39:27]
  wire  _T_398; // @[LZD.scala 39:25]
  wire [1:0] _T_399; // @[Cat.scala 29:58]
  wire [1:0] _T_400; // @[LZD.scala 44:32]
  wire  _T_401; // @[LZD.scala 39:14]
  wire  _T_402; // @[LZD.scala 39:21]
  wire  _T_403; // @[LZD.scala 39:30]
  wire  _T_404; // @[LZD.scala 39:27]
  wire  _T_405; // @[LZD.scala 39:25]
  wire [1:0] _T_406; // @[Cat.scala 29:58]
  wire  _T_407; // @[Shift.scala 12:21]
  wire  _T_408; // @[Shift.scala 12:21]
  wire  _T_409; // @[LZD.scala 49:16]
  wire  _T_410; // @[LZD.scala 49:27]
  wire  _T_411; // @[LZD.scala 49:25]
  wire  _T_412; // @[LZD.scala 49:47]
  wire  _T_413; // @[LZD.scala 49:59]
  wire  _T_414; // @[LZD.scala 49:35]
  wire [2:0] _T_416; // @[Cat.scala 29:58]
  wire  _T_417; // @[Shift.scala 12:21]
  wire  _T_418; // @[Shift.scala 12:21]
  wire  _T_419; // @[LZD.scala 49:16]
  wire  _T_420; // @[LZD.scala 49:27]
  wire  _T_421; // @[LZD.scala 49:25]
  wire [1:0] _T_422; // @[LZD.scala 49:47]
  wire [1:0] _T_423; // @[LZD.scala 49:59]
  wire [1:0] _T_424; // @[LZD.scala 49:35]
  wire [3:0] _T_426; // @[Cat.scala 29:58]
  wire  _T_427; // @[Shift.scala 12:21]
  wire  _T_428; // @[Shift.scala 12:21]
  wire  _T_429; // @[LZD.scala 49:16]
  wire  _T_430; // @[LZD.scala 49:27]
  wire  _T_431; // @[LZD.scala 49:25]
  wire [2:0] _T_432; // @[LZD.scala 49:47]
  wire [2:0] _T_433; // @[LZD.scala 49:59]
  wire [2:0] _T_434; // @[LZD.scala 49:35]
  wire [4:0] _T_436; // @[Cat.scala 29:58]
  wire [10:0] _T_437; // @[LZD.scala 44:32]
  wire [7:0] _T_438; // @[LZD.scala 43:32]
  wire [3:0] _T_439; // @[LZD.scala 43:32]
  wire [1:0] _T_440; // @[LZD.scala 43:32]
  wire  _T_441; // @[LZD.scala 39:14]
  wire  _T_442; // @[LZD.scala 39:21]
  wire  _T_443; // @[LZD.scala 39:30]
  wire  _T_444; // @[LZD.scala 39:27]
  wire  _T_445; // @[LZD.scala 39:25]
  wire [1:0] _T_446; // @[Cat.scala 29:58]
  wire [1:0] _T_447; // @[LZD.scala 44:32]
  wire  _T_448; // @[LZD.scala 39:14]
  wire  _T_449; // @[LZD.scala 39:21]
  wire  _T_450; // @[LZD.scala 39:30]
  wire  _T_451; // @[LZD.scala 39:27]
  wire  _T_452; // @[LZD.scala 39:25]
  wire [1:0] _T_453; // @[Cat.scala 29:58]
  wire  _T_454; // @[Shift.scala 12:21]
  wire  _T_455; // @[Shift.scala 12:21]
  wire  _T_456; // @[LZD.scala 49:16]
  wire  _T_457; // @[LZD.scala 49:27]
  wire  _T_458; // @[LZD.scala 49:25]
  wire  _T_459; // @[LZD.scala 49:47]
  wire  _T_460; // @[LZD.scala 49:59]
  wire  _T_461; // @[LZD.scala 49:35]
  wire [2:0] _T_463; // @[Cat.scala 29:58]
  wire [3:0] _T_464; // @[LZD.scala 44:32]
  wire [1:0] _T_465; // @[LZD.scala 43:32]
  wire  _T_466; // @[LZD.scala 39:14]
  wire  _T_467; // @[LZD.scala 39:21]
  wire  _T_468; // @[LZD.scala 39:30]
  wire  _T_469; // @[LZD.scala 39:27]
  wire  _T_470; // @[LZD.scala 39:25]
  wire [1:0] _T_471; // @[Cat.scala 29:58]
  wire [1:0] _T_472; // @[LZD.scala 44:32]
  wire  _T_473; // @[LZD.scala 39:14]
  wire  _T_474; // @[LZD.scala 39:21]
  wire  _T_475; // @[LZD.scala 39:30]
  wire  _T_476; // @[LZD.scala 39:27]
  wire  _T_477; // @[LZD.scala 39:25]
  wire [1:0] _T_478; // @[Cat.scala 29:58]
  wire  _T_479; // @[Shift.scala 12:21]
  wire  _T_480; // @[Shift.scala 12:21]
  wire  _T_481; // @[LZD.scala 49:16]
  wire  _T_482; // @[LZD.scala 49:27]
  wire  _T_483; // @[LZD.scala 49:25]
  wire  _T_484; // @[LZD.scala 49:47]
  wire  _T_485; // @[LZD.scala 49:59]
  wire  _T_486; // @[LZD.scala 49:35]
  wire [2:0] _T_488; // @[Cat.scala 29:58]
  wire  _T_489; // @[Shift.scala 12:21]
  wire  _T_490; // @[Shift.scala 12:21]
  wire  _T_491; // @[LZD.scala 49:16]
  wire  _T_492; // @[LZD.scala 49:27]
  wire  _T_493; // @[LZD.scala 49:25]
  wire [1:0] _T_494; // @[LZD.scala 49:47]
  wire [1:0] _T_495; // @[LZD.scala 49:59]
  wire [1:0] _T_496; // @[LZD.scala 49:35]
  wire [3:0] _T_498; // @[Cat.scala 29:58]
  wire [2:0] _T_499; // @[LZD.scala 44:32]
  wire [1:0] _T_500; // @[LZD.scala 43:32]
  wire  _T_501; // @[LZD.scala 39:14]
  wire  _T_502; // @[LZD.scala 39:21]
  wire  _T_503; // @[LZD.scala 39:30]
  wire  _T_504; // @[LZD.scala 39:27]
  wire  _T_505; // @[LZD.scala 39:25]
  wire [1:0] _T_506; // @[Cat.scala 29:58]
  wire  _T_507; // @[LZD.scala 44:32]
  wire  _T_509; // @[Shift.scala 12:21]
  wire  _T_511; // @[LZD.scala 55:32]
  wire  _T_512; // @[LZD.scala 55:20]
  wire  _T_514; // @[Shift.scala 12:21]
  wire [2:0] _T_516; // @[Cat.scala 29:58]
  wire [2:0] _T_517; // @[LZD.scala 55:32]
  wire [2:0] _T_518; // @[LZD.scala 55:20]
  wire [3:0] _T_519; // @[Cat.scala 29:58]
  wire  _T_520; // @[Shift.scala 12:21]
  wire [3:0] _T_522; // @[LZD.scala 55:32]
  wire [3:0] _T_523; // @[LZD.scala 55:20]
  wire [4:0] _T_524; // @[Cat.scala 29:58]
  wire [4:0] _T_525; // @[convert.scala 21:22]
  wire [25:0] _T_526; // @[convert.scala 22:36]
  wire  _T_527; // @[Shift.scala 16:24]
  wire  _T_529; // @[Shift.scala 12:21]
  wire [9:0] _T_530; // @[Shift.scala 64:52]
  wire [25:0] _T_532; // @[Cat.scala 29:58]
  wire [25:0] _T_533; // @[Shift.scala 64:27]
  wire [3:0] _T_534; // @[Shift.scala 66:70]
  wire  _T_535; // @[Shift.scala 12:21]
  wire [17:0] _T_536; // @[Shift.scala 64:52]
  wire [25:0] _T_538; // @[Cat.scala 29:58]
  wire [25:0] _T_539; // @[Shift.scala 64:27]
  wire [2:0] _T_540; // @[Shift.scala 66:70]
  wire  _T_541; // @[Shift.scala 12:21]
  wire [21:0] _T_542; // @[Shift.scala 64:52]
  wire [25:0] _T_544; // @[Cat.scala 29:58]
  wire [25:0] _T_545; // @[Shift.scala 64:27]
  wire [1:0] _T_546; // @[Shift.scala 66:70]
  wire  _T_547; // @[Shift.scala 12:21]
  wire [23:0] _T_548; // @[Shift.scala 64:52]
  wire [25:0] _T_550; // @[Cat.scala 29:58]
  wire [25:0] _T_551; // @[Shift.scala 64:27]
  wire  _T_552; // @[Shift.scala 66:70]
  wire [24:0] _T_554; // @[Shift.scala 64:52]
  wire [25:0] _T_555; // @[Cat.scala 29:58]
  wire [25:0] _T_556; // @[Shift.scala 64:27]
  wire [25:0] _T_557; // @[Shift.scala 16:10]
  wire [2:0] _T_558; // @[convert.scala 23:34]
  wire [22:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_560; // @[convert.scala 25:26]
  wire [4:0] _T_562; // @[convert.scala 25:42]
  wire [2:0] _T_565; // @[convert.scala 26:67]
  wire [2:0] _T_566; // @[convert.scala 26:51]
  wire [8:0] _T_567; // @[Cat.scala 29:58]
  wire [27:0] _T_569; // @[convert.scala 29:56]
  wire  _T_570; // @[convert.scala 29:60]
  wire  _T_571; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_574; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [8:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_583; // @[convert.scala 18:24]
  wire  _T_584; // @[convert.scala 18:40]
  wire  _T_585; // @[convert.scala 18:36]
  wire [26:0] _T_586; // @[convert.scala 19:24]
  wire [26:0] _T_587; // @[convert.scala 19:43]
  wire [26:0] _T_588; // @[convert.scala 19:39]
  wire [15:0] _T_589; // @[LZD.scala 43:32]
  wire [7:0] _T_590; // @[LZD.scala 43:32]
  wire [3:0] _T_591; // @[LZD.scala 43:32]
  wire [1:0] _T_592; // @[LZD.scala 43:32]
  wire  _T_593; // @[LZD.scala 39:14]
  wire  _T_594; // @[LZD.scala 39:21]
  wire  _T_595; // @[LZD.scala 39:30]
  wire  _T_596; // @[LZD.scala 39:27]
  wire  _T_597; // @[LZD.scala 39:25]
  wire [1:0] _T_598; // @[Cat.scala 29:58]
  wire [1:0] _T_599; // @[LZD.scala 44:32]
  wire  _T_600; // @[LZD.scala 39:14]
  wire  _T_601; // @[LZD.scala 39:21]
  wire  _T_602; // @[LZD.scala 39:30]
  wire  _T_603; // @[LZD.scala 39:27]
  wire  _T_604; // @[LZD.scala 39:25]
  wire [1:0] _T_605; // @[Cat.scala 29:58]
  wire  _T_606; // @[Shift.scala 12:21]
  wire  _T_607; // @[Shift.scala 12:21]
  wire  _T_608; // @[LZD.scala 49:16]
  wire  _T_609; // @[LZD.scala 49:27]
  wire  _T_610; // @[LZD.scala 49:25]
  wire  _T_611; // @[LZD.scala 49:47]
  wire  _T_612; // @[LZD.scala 49:59]
  wire  _T_613; // @[LZD.scala 49:35]
  wire [2:0] _T_615; // @[Cat.scala 29:58]
  wire [3:0] _T_616; // @[LZD.scala 44:32]
  wire [1:0] _T_617; // @[LZD.scala 43:32]
  wire  _T_618; // @[LZD.scala 39:14]
  wire  _T_619; // @[LZD.scala 39:21]
  wire  _T_620; // @[LZD.scala 39:30]
  wire  _T_621; // @[LZD.scala 39:27]
  wire  _T_622; // @[LZD.scala 39:25]
  wire [1:0] _T_623; // @[Cat.scala 29:58]
  wire [1:0] _T_624; // @[LZD.scala 44:32]
  wire  _T_625; // @[LZD.scala 39:14]
  wire  _T_626; // @[LZD.scala 39:21]
  wire  _T_627; // @[LZD.scala 39:30]
  wire  _T_628; // @[LZD.scala 39:27]
  wire  _T_629; // @[LZD.scala 39:25]
  wire [1:0] _T_630; // @[Cat.scala 29:58]
  wire  _T_631; // @[Shift.scala 12:21]
  wire  _T_632; // @[Shift.scala 12:21]
  wire  _T_633; // @[LZD.scala 49:16]
  wire  _T_634; // @[LZD.scala 49:27]
  wire  _T_635; // @[LZD.scala 49:25]
  wire  _T_636; // @[LZD.scala 49:47]
  wire  _T_637; // @[LZD.scala 49:59]
  wire  _T_638; // @[LZD.scala 49:35]
  wire [2:0] _T_640; // @[Cat.scala 29:58]
  wire  _T_641; // @[Shift.scala 12:21]
  wire  _T_642; // @[Shift.scala 12:21]
  wire  _T_643; // @[LZD.scala 49:16]
  wire  _T_644; // @[LZD.scala 49:27]
  wire  _T_645; // @[LZD.scala 49:25]
  wire [1:0] _T_646; // @[LZD.scala 49:47]
  wire [1:0] _T_647; // @[LZD.scala 49:59]
  wire [1:0] _T_648; // @[LZD.scala 49:35]
  wire [3:0] _T_650; // @[Cat.scala 29:58]
  wire [7:0] _T_651; // @[LZD.scala 44:32]
  wire [3:0] _T_652; // @[LZD.scala 43:32]
  wire [1:0] _T_653; // @[LZD.scala 43:32]
  wire  _T_654; // @[LZD.scala 39:14]
  wire  _T_655; // @[LZD.scala 39:21]
  wire  _T_656; // @[LZD.scala 39:30]
  wire  _T_657; // @[LZD.scala 39:27]
  wire  _T_658; // @[LZD.scala 39:25]
  wire [1:0] _T_659; // @[Cat.scala 29:58]
  wire [1:0] _T_660; // @[LZD.scala 44:32]
  wire  _T_661; // @[LZD.scala 39:14]
  wire  _T_662; // @[LZD.scala 39:21]
  wire  _T_663; // @[LZD.scala 39:30]
  wire  _T_664; // @[LZD.scala 39:27]
  wire  _T_665; // @[LZD.scala 39:25]
  wire [1:0] _T_666; // @[Cat.scala 29:58]
  wire  _T_667; // @[Shift.scala 12:21]
  wire  _T_668; // @[Shift.scala 12:21]
  wire  _T_669; // @[LZD.scala 49:16]
  wire  _T_670; // @[LZD.scala 49:27]
  wire  _T_671; // @[LZD.scala 49:25]
  wire  _T_672; // @[LZD.scala 49:47]
  wire  _T_673; // @[LZD.scala 49:59]
  wire  _T_674; // @[LZD.scala 49:35]
  wire [2:0] _T_676; // @[Cat.scala 29:58]
  wire [3:0] _T_677; // @[LZD.scala 44:32]
  wire [1:0] _T_678; // @[LZD.scala 43:32]
  wire  _T_679; // @[LZD.scala 39:14]
  wire  _T_680; // @[LZD.scala 39:21]
  wire  _T_681; // @[LZD.scala 39:30]
  wire  _T_682; // @[LZD.scala 39:27]
  wire  _T_683; // @[LZD.scala 39:25]
  wire [1:0] _T_684; // @[Cat.scala 29:58]
  wire [1:0] _T_685; // @[LZD.scala 44:32]
  wire  _T_686; // @[LZD.scala 39:14]
  wire  _T_687; // @[LZD.scala 39:21]
  wire  _T_688; // @[LZD.scala 39:30]
  wire  _T_689; // @[LZD.scala 39:27]
  wire  _T_690; // @[LZD.scala 39:25]
  wire [1:0] _T_691; // @[Cat.scala 29:58]
  wire  _T_692; // @[Shift.scala 12:21]
  wire  _T_693; // @[Shift.scala 12:21]
  wire  _T_694; // @[LZD.scala 49:16]
  wire  _T_695; // @[LZD.scala 49:27]
  wire  _T_696; // @[LZD.scala 49:25]
  wire  _T_697; // @[LZD.scala 49:47]
  wire  _T_698; // @[LZD.scala 49:59]
  wire  _T_699; // @[LZD.scala 49:35]
  wire [2:0] _T_701; // @[Cat.scala 29:58]
  wire  _T_702; // @[Shift.scala 12:21]
  wire  _T_703; // @[Shift.scala 12:21]
  wire  _T_704; // @[LZD.scala 49:16]
  wire  _T_705; // @[LZD.scala 49:27]
  wire  _T_706; // @[LZD.scala 49:25]
  wire [1:0] _T_707; // @[LZD.scala 49:47]
  wire [1:0] _T_708; // @[LZD.scala 49:59]
  wire [1:0] _T_709; // @[LZD.scala 49:35]
  wire [3:0] _T_711; // @[Cat.scala 29:58]
  wire  _T_712; // @[Shift.scala 12:21]
  wire  _T_713; // @[Shift.scala 12:21]
  wire  _T_714; // @[LZD.scala 49:16]
  wire  _T_715; // @[LZD.scala 49:27]
  wire  _T_716; // @[LZD.scala 49:25]
  wire [2:0] _T_717; // @[LZD.scala 49:47]
  wire [2:0] _T_718; // @[LZD.scala 49:59]
  wire [2:0] _T_719; // @[LZD.scala 49:35]
  wire [4:0] _T_721; // @[Cat.scala 29:58]
  wire [10:0] _T_722; // @[LZD.scala 44:32]
  wire [7:0] _T_723; // @[LZD.scala 43:32]
  wire [3:0] _T_724; // @[LZD.scala 43:32]
  wire [1:0] _T_725; // @[LZD.scala 43:32]
  wire  _T_726; // @[LZD.scala 39:14]
  wire  _T_727; // @[LZD.scala 39:21]
  wire  _T_728; // @[LZD.scala 39:30]
  wire  _T_729; // @[LZD.scala 39:27]
  wire  _T_730; // @[LZD.scala 39:25]
  wire [1:0] _T_731; // @[Cat.scala 29:58]
  wire [1:0] _T_732; // @[LZD.scala 44:32]
  wire  _T_733; // @[LZD.scala 39:14]
  wire  _T_734; // @[LZD.scala 39:21]
  wire  _T_735; // @[LZD.scala 39:30]
  wire  _T_736; // @[LZD.scala 39:27]
  wire  _T_737; // @[LZD.scala 39:25]
  wire [1:0] _T_738; // @[Cat.scala 29:58]
  wire  _T_739; // @[Shift.scala 12:21]
  wire  _T_740; // @[Shift.scala 12:21]
  wire  _T_741; // @[LZD.scala 49:16]
  wire  _T_742; // @[LZD.scala 49:27]
  wire  _T_743; // @[LZD.scala 49:25]
  wire  _T_744; // @[LZD.scala 49:47]
  wire  _T_745; // @[LZD.scala 49:59]
  wire  _T_746; // @[LZD.scala 49:35]
  wire [2:0] _T_748; // @[Cat.scala 29:58]
  wire [3:0] _T_749; // @[LZD.scala 44:32]
  wire [1:0] _T_750; // @[LZD.scala 43:32]
  wire  _T_751; // @[LZD.scala 39:14]
  wire  _T_752; // @[LZD.scala 39:21]
  wire  _T_753; // @[LZD.scala 39:30]
  wire  _T_754; // @[LZD.scala 39:27]
  wire  _T_755; // @[LZD.scala 39:25]
  wire [1:0] _T_756; // @[Cat.scala 29:58]
  wire [1:0] _T_757; // @[LZD.scala 44:32]
  wire  _T_758; // @[LZD.scala 39:14]
  wire  _T_759; // @[LZD.scala 39:21]
  wire  _T_760; // @[LZD.scala 39:30]
  wire  _T_761; // @[LZD.scala 39:27]
  wire  _T_762; // @[LZD.scala 39:25]
  wire [1:0] _T_763; // @[Cat.scala 29:58]
  wire  _T_764; // @[Shift.scala 12:21]
  wire  _T_765; // @[Shift.scala 12:21]
  wire  _T_766; // @[LZD.scala 49:16]
  wire  _T_767; // @[LZD.scala 49:27]
  wire  _T_768; // @[LZD.scala 49:25]
  wire  _T_769; // @[LZD.scala 49:47]
  wire  _T_770; // @[LZD.scala 49:59]
  wire  _T_771; // @[LZD.scala 49:35]
  wire [2:0] _T_773; // @[Cat.scala 29:58]
  wire  _T_774; // @[Shift.scala 12:21]
  wire  _T_775; // @[Shift.scala 12:21]
  wire  _T_776; // @[LZD.scala 49:16]
  wire  _T_777; // @[LZD.scala 49:27]
  wire  _T_778; // @[LZD.scala 49:25]
  wire [1:0] _T_779; // @[LZD.scala 49:47]
  wire [1:0] _T_780; // @[LZD.scala 49:59]
  wire [1:0] _T_781; // @[LZD.scala 49:35]
  wire [3:0] _T_783; // @[Cat.scala 29:58]
  wire [2:0] _T_784; // @[LZD.scala 44:32]
  wire [1:0] _T_785; // @[LZD.scala 43:32]
  wire  _T_786; // @[LZD.scala 39:14]
  wire  _T_787; // @[LZD.scala 39:21]
  wire  _T_788; // @[LZD.scala 39:30]
  wire  _T_789; // @[LZD.scala 39:27]
  wire  _T_790; // @[LZD.scala 39:25]
  wire [1:0] _T_791; // @[Cat.scala 29:58]
  wire  _T_792; // @[LZD.scala 44:32]
  wire  _T_794; // @[Shift.scala 12:21]
  wire  _T_796; // @[LZD.scala 55:32]
  wire  _T_797; // @[LZD.scala 55:20]
  wire  _T_799; // @[Shift.scala 12:21]
  wire [2:0] _T_801; // @[Cat.scala 29:58]
  wire [2:0] _T_802; // @[LZD.scala 55:32]
  wire [2:0] _T_803; // @[LZD.scala 55:20]
  wire [3:0] _T_804; // @[Cat.scala 29:58]
  wire  _T_805; // @[Shift.scala 12:21]
  wire [3:0] _T_807; // @[LZD.scala 55:32]
  wire [3:0] _T_808; // @[LZD.scala 55:20]
  wire [4:0] _T_809; // @[Cat.scala 29:58]
  wire [4:0] _T_810; // @[convert.scala 21:22]
  wire [25:0] _T_811; // @[convert.scala 22:36]
  wire  _T_812; // @[Shift.scala 16:24]
  wire  _T_814; // @[Shift.scala 12:21]
  wire [9:0] _T_815; // @[Shift.scala 64:52]
  wire [25:0] _T_817; // @[Cat.scala 29:58]
  wire [25:0] _T_818; // @[Shift.scala 64:27]
  wire [3:0] _T_819; // @[Shift.scala 66:70]
  wire  _T_820; // @[Shift.scala 12:21]
  wire [17:0] _T_821; // @[Shift.scala 64:52]
  wire [25:0] _T_823; // @[Cat.scala 29:58]
  wire [25:0] _T_824; // @[Shift.scala 64:27]
  wire [2:0] _T_825; // @[Shift.scala 66:70]
  wire  _T_826; // @[Shift.scala 12:21]
  wire [21:0] _T_827; // @[Shift.scala 64:52]
  wire [25:0] _T_829; // @[Cat.scala 29:58]
  wire [25:0] _T_830; // @[Shift.scala 64:27]
  wire [1:0] _T_831; // @[Shift.scala 66:70]
  wire  _T_832; // @[Shift.scala 12:21]
  wire [23:0] _T_833; // @[Shift.scala 64:52]
  wire [25:0] _T_835; // @[Cat.scala 29:58]
  wire [25:0] _T_836; // @[Shift.scala 64:27]
  wire  _T_837; // @[Shift.scala 66:70]
  wire [24:0] _T_839; // @[Shift.scala 64:52]
  wire [25:0] _T_840; // @[Cat.scala 29:58]
  wire [25:0] _T_841; // @[Shift.scala 64:27]
  wire [25:0] _T_842; // @[Shift.scala 16:10]
  wire [2:0] _T_843; // @[convert.scala 23:34]
  wire [22:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_845; // @[convert.scala 25:26]
  wire [4:0] _T_847; // @[convert.scala 25:42]
  wire [2:0] _T_850; // @[convert.scala 26:67]
  wire [2:0] _T_851; // @[convert.scala 26:51]
  wire [8:0] _T_852; // @[Cat.scala 29:58]
  wire [27:0] _T_854; // @[convert.scala 29:56]
  wire  _T_855; // @[convert.scala 29:60]
  wire  _T_856; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_859; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [8:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_867; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_868; // @[PositFMA.scala 59:34]
  wire  _T_869; // @[PositFMA.scala 59:47]
  wire  _T_870; // @[PositFMA.scala 59:45]
  wire [24:0] _T_872; // @[Cat.scala 29:58]
  wire [24:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_873; // @[PositFMA.scala 60:34]
  wire  _T_874; // @[PositFMA.scala 60:47]
  wire  _T_875; // @[PositFMA.scala 60:45]
  wire [24:0] _T_877; // @[Cat.scala 29:58]
  wire [24:0] sigB; // @[PositFMA.scala 60:76]
  wire [49:0] _T_878; // @[PositFMA.scala 61:25]
  wire [49:0] sigP; // @[PositFMA.scala 61:33]
  wire [46:0] _T_879; // @[PositFMA.scala 62:29]
  wire  _T_880; // @[PositFMA.scala 62:33]
  wire  eqTwo; // @[PositFMA.scala 62:19]
  wire  _T_881; // @[PositFMA.scala 64:29]
  wire  _T_882; // @[PositFMA.scala 64:56]
  wire  _T_883; // @[PositFMA.scala 64:51]
  wire  _T_884; // @[PositFMA.scala 64:49]
  wire  eqFour; // @[PositFMA.scala 64:76]
  wire  _T_885; // @[PositFMA.scala 66:23]
  wire  geTwo; // @[PositFMA.scala 66:43]
  wire [1:0] _T_887; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 67:38]
  wire  mulSign; // @[PositFMA.scala 68:28]
  wire [9:0] _T_888; // @[PositFMA.scala 70:30]
  wire [9:0] _GEN_12; // @[PositFMA.scala 70:44]
  wire [9:0] _T_890; // @[PositFMA.scala 70:44]
  wire [9:0] mulScale; // @[PositFMA.scala 70:44]
  wire [47:0] _T_891; // @[PositFMA.scala 73:29]
  wire [46:0] _T_892; // @[PositFMA.scala 74:29]
  wire [47:0] _T_893; // @[PositFMA.scala 74:48]
  wire [47:0] mulSigTmp; // @[PositFMA.scala 71:22]
  wire  _T_895; // @[PositFMA.scala 78:39]
  wire  _T_896; // @[PositFMA.scala 78:43]
  wire [46:0] _T_897; // @[PositFMA.scala 79:39]
  wire [48:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [48:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [63:0] _RAND_1;
  reg [22:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [9:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [8:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_923; // @[PositFMA.scala 108:29]
  wire  _T_924; // @[PositFMA.scala 108:47]
  wire  _T_925; // @[PositFMA.scala 108:45]
  wire [48:0] extAddSig; // @[Cat.scala 29:58]
  wire [9:0] _GEN_13; // @[PositFMA.scala 112:39]
  wire  mulGreater; // @[PositFMA.scala 112:39]
  wire [9:0] greaterScale; // @[PositFMA.scala 113:26]
  wire [9:0] smallerScale; // @[PositFMA.scala 114:26]
  wire [9:0] _T_929; // @[PositFMA.scala 115:36]
  wire [9:0] scaleDiff; // @[PositFMA.scala 115:36]
  wire [48:0] greaterSig; // @[PositFMA.scala 116:26]
  wire [48:0] smallerSigTmp; // @[PositFMA.scala 117:26]
  wire [9:0] _T_930; // @[PositFMA.scala 118:69]
  wire  _T_931; // @[Shift.scala 39:24]
  wire [5:0] _T_932; // @[Shift.scala 40:44]
  wire [16:0] _T_933; // @[Shift.scala 90:30]
  wire [31:0] _T_934; // @[Shift.scala 90:48]
  wire  _T_935; // @[Shift.scala 90:57]
  wire [16:0] _GEN_14; // @[Shift.scala 90:39]
  wire [16:0] _T_936; // @[Shift.scala 90:39]
  wire  _T_937; // @[Shift.scala 12:21]
  wire  _T_938; // @[Shift.scala 12:21]
  wire [31:0] _T_940; // @[Bitwise.scala 71:12]
  wire [48:0] _T_941; // @[Cat.scala 29:58]
  wire [48:0] _T_942; // @[Shift.scala 91:22]
  wire [4:0] _T_943; // @[Shift.scala 92:77]
  wire [32:0] _T_944; // @[Shift.scala 90:30]
  wire [15:0] _T_945; // @[Shift.scala 90:48]
  wire  _T_946; // @[Shift.scala 90:57]
  wire [32:0] _GEN_15; // @[Shift.scala 90:39]
  wire [32:0] _T_947; // @[Shift.scala 90:39]
  wire  _T_948; // @[Shift.scala 12:21]
  wire  _T_949; // @[Shift.scala 12:21]
  wire [15:0] _T_951; // @[Bitwise.scala 71:12]
  wire [48:0] _T_952; // @[Cat.scala 29:58]
  wire [48:0] _T_953; // @[Shift.scala 91:22]
  wire [3:0] _T_954; // @[Shift.scala 92:77]
  wire [40:0] _T_955; // @[Shift.scala 90:30]
  wire [7:0] _T_956; // @[Shift.scala 90:48]
  wire  _T_957; // @[Shift.scala 90:57]
  wire [40:0] _GEN_16; // @[Shift.scala 90:39]
  wire [40:0] _T_958; // @[Shift.scala 90:39]
  wire  _T_959; // @[Shift.scala 12:21]
  wire  _T_960; // @[Shift.scala 12:21]
  wire [7:0] _T_962; // @[Bitwise.scala 71:12]
  wire [48:0] _T_963; // @[Cat.scala 29:58]
  wire [48:0] _T_964; // @[Shift.scala 91:22]
  wire [2:0] _T_965; // @[Shift.scala 92:77]
  wire [44:0] _T_966; // @[Shift.scala 90:30]
  wire [3:0] _T_967; // @[Shift.scala 90:48]
  wire  _T_968; // @[Shift.scala 90:57]
  wire [44:0] _GEN_17; // @[Shift.scala 90:39]
  wire [44:0] _T_969; // @[Shift.scala 90:39]
  wire  _T_970; // @[Shift.scala 12:21]
  wire  _T_971; // @[Shift.scala 12:21]
  wire [3:0] _T_973; // @[Bitwise.scala 71:12]
  wire [48:0] _T_974; // @[Cat.scala 29:58]
  wire [48:0] _T_975; // @[Shift.scala 91:22]
  wire [1:0] _T_976; // @[Shift.scala 92:77]
  wire [46:0] _T_977; // @[Shift.scala 90:30]
  wire [1:0] _T_978; // @[Shift.scala 90:48]
  wire  _T_979; // @[Shift.scala 90:57]
  wire [46:0] _GEN_18; // @[Shift.scala 90:39]
  wire [46:0] _T_980; // @[Shift.scala 90:39]
  wire  _T_981; // @[Shift.scala 12:21]
  wire  _T_982; // @[Shift.scala 12:21]
  wire [1:0] _T_984; // @[Bitwise.scala 71:12]
  wire [48:0] _T_985; // @[Cat.scala 29:58]
  wire [48:0] _T_986; // @[Shift.scala 91:22]
  wire  _T_987; // @[Shift.scala 92:77]
  wire [47:0] _T_988; // @[Shift.scala 90:30]
  wire  _T_989; // @[Shift.scala 90:48]
  wire [47:0] _GEN_19; // @[Shift.scala 90:39]
  wire [47:0] _T_991; // @[Shift.scala 90:39]
  wire  _T_993; // @[Shift.scala 12:21]
  wire [48:0] _T_994; // @[Cat.scala 29:58]
  wire [48:0] _T_995; // @[Shift.scala 91:22]
  wire [48:0] _T_998; // @[Bitwise.scala 71:12]
  wire [48:0] smallerSig; // @[Shift.scala 39:10]
  wire [49:0] rawSumSig; // @[PositFMA.scala 119:34]
  wire  _T_999; // @[PositFMA.scala 120:42]
  wire  _T_1000; // @[PositFMA.scala 120:46]
  wire  _T_1001; // @[PositFMA.scala 120:79]
  wire  sumSign; // @[PositFMA.scala 120:63]
  wire [48:0] _T_1003; // @[PositFMA.scala 121:50]
  wire [49:0] signSumSig; // @[Cat.scala 29:58]
  wire [48:0] _T_1004; // @[PositFMA.scala 125:33]
  wire [48:0] _T_1005; // @[PositFMA.scala 125:68]
  wire [48:0] sumXor; // @[PositFMA.scala 125:51]
  wire [31:0] _T_1006; // @[LZD.scala 43:32]
  wire [15:0] _T_1007; // @[LZD.scala 43:32]
  wire [7:0] _T_1008; // @[LZD.scala 43:32]
  wire [3:0] _T_1009; // @[LZD.scala 43:32]
  wire [1:0] _T_1010; // @[LZD.scala 43:32]
  wire  _T_1011; // @[LZD.scala 39:14]
  wire  _T_1012; // @[LZD.scala 39:21]
  wire  _T_1013; // @[LZD.scala 39:30]
  wire  _T_1014; // @[LZD.scala 39:27]
  wire  _T_1015; // @[LZD.scala 39:25]
  wire [1:0] _T_1016; // @[Cat.scala 29:58]
  wire [1:0] _T_1017; // @[LZD.scala 44:32]
  wire  _T_1018; // @[LZD.scala 39:14]
  wire  _T_1019; // @[LZD.scala 39:21]
  wire  _T_1020; // @[LZD.scala 39:30]
  wire  _T_1021; // @[LZD.scala 39:27]
  wire  _T_1022; // @[LZD.scala 39:25]
  wire [1:0] _T_1023; // @[Cat.scala 29:58]
  wire  _T_1024; // @[Shift.scala 12:21]
  wire  _T_1025; // @[Shift.scala 12:21]
  wire  _T_1026; // @[LZD.scala 49:16]
  wire  _T_1027; // @[LZD.scala 49:27]
  wire  _T_1028; // @[LZD.scala 49:25]
  wire  _T_1029; // @[LZD.scala 49:47]
  wire  _T_1030; // @[LZD.scala 49:59]
  wire  _T_1031; // @[LZD.scala 49:35]
  wire [2:0] _T_1033; // @[Cat.scala 29:58]
  wire [3:0] _T_1034; // @[LZD.scala 44:32]
  wire [1:0] _T_1035; // @[LZD.scala 43:32]
  wire  _T_1036; // @[LZD.scala 39:14]
  wire  _T_1037; // @[LZD.scala 39:21]
  wire  _T_1038; // @[LZD.scala 39:30]
  wire  _T_1039; // @[LZD.scala 39:27]
  wire  _T_1040; // @[LZD.scala 39:25]
  wire [1:0] _T_1041; // @[Cat.scala 29:58]
  wire [1:0] _T_1042; // @[LZD.scala 44:32]
  wire  _T_1043; // @[LZD.scala 39:14]
  wire  _T_1044; // @[LZD.scala 39:21]
  wire  _T_1045; // @[LZD.scala 39:30]
  wire  _T_1046; // @[LZD.scala 39:27]
  wire  _T_1047; // @[LZD.scala 39:25]
  wire [1:0] _T_1048; // @[Cat.scala 29:58]
  wire  _T_1049; // @[Shift.scala 12:21]
  wire  _T_1050; // @[Shift.scala 12:21]
  wire  _T_1051; // @[LZD.scala 49:16]
  wire  _T_1052; // @[LZD.scala 49:27]
  wire  _T_1053; // @[LZD.scala 49:25]
  wire  _T_1054; // @[LZD.scala 49:47]
  wire  _T_1055; // @[LZD.scala 49:59]
  wire  _T_1056; // @[LZD.scala 49:35]
  wire [2:0] _T_1058; // @[Cat.scala 29:58]
  wire  _T_1059; // @[Shift.scala 12:21]
  wire  _T_1060; // @[Shift.scala 12:21]
  wire  _T_1061; // @[LZD.scala 49:16]
  wire  _T_1062; // @[LZD.scala 49:27]
  wire  _T_1063; // @[LZD.scala 49:25]
  wire [1:0] _T_1064; // @[LZD.scala 49:47]
  wire [1:0] _T_1065; // @[LZD.scala 49:59]
  wire [1:0] _T_1066; // @[LZD.scala 49:35]
  wire [3:0] _T_1068; // @[Cat.scala 29:58]
  wire [7:0] _T_1069; // @[LZD.scala 44:32]
  wire [3:0] _T_1070; // @[LZD.scala 43:32]
  wire [1:0] _T_1071; // @[LZD.scala 43:32]
  wire  _T_1072; // @[LZD.scala 39:14]
  wire  _T_1073; // @[LZD.scala 39:21]
  wire  _T_1074; // @[LZD.scala 39:30]
  wire  _T_1075; // @[LZD.scala 39:27]
  wire  _T_1076; // @[LZD.scala 39:25]
  wire [1:0] _T_1077; // @[Cat.scala 29:58]
  wire [1:0] _T_1078; // @[LZD.scala 44:32]
  wire  _T_1079; // @[LZD.scala 39:14]
  wire  _T_1080; // @[LZD.scala 39:21]
  wire  _T_1081; // @[LZD.scala 39:30]
  wire  _T_1082; // @[LZD.scala 39:27]
  wire  _T_1083; // @[LZD.scala 39:25]
  wire [1:0] _T_1084; // @[Cat.scala 29:58]
  wire  _T_1085; // @[Shift.scala 12:21]
  wire  _T_1086; // @[Shift.scala 12:21]
  wire  _T_1087; // @[LZD.scala 49:16]
  wire  _T_1088; // @[LZD.scala 49:27]
  wire  _T_1089; // @[LZD.scala 49:25]
  wire  _T_1090; // @[LZD.scala 49:47]
  wire  _T_1091; // @[LZD.scala 49:59]
  wire  _T_1092; // @[LZD.scala 49:35]
  wire [2:0] _T_1094; // @[Cat.scala 29:58]
  wire [3:0] _T_1095; // @[LZD.scala 44:32]
  wire [1:0] _T_1096; // @[LZD.scala 43:32]
  wire  _T_1097; // @[LZD.scala 39:14]
  wire  _T_1098; // @[LZD.scala 39:21]
  wire  _T_1099; // @[LZD.scala 39:30]
  wire  _T_1100; // @[LZD.scala 39:27]
  wire  _T_1101; // @[LZD.scala 39:25]
  wire [1:0] _T_1102; // @[Cat.scala 29:58]
  wire [1:0] _T_1103; // @[LZD.scala 44:32]
  wire  _T_1104; // @[LZD.scala 39:14]
  wire  _T_1105; // @[LZD.scala 39:21]
  wire  _T_1106; // @[LZD.scala 39:30]
  wire  _T_1107; // @[LZD.scala 39:27]
  wire  _T_1108; // @[LZD.scala 39:25]
  wire [1:0] _T_1109; // @[Cat.scala 29:58]
  wire  _T_1110; // @[Shift.scala 12:21]
  wire  _T_1111; // @[Shift.scala 12:21]
  wire  _T_1112; // @[LZD.scala 49:16]
  wire  _T_1113; // @[LZD.scala 49:27]
  wire  _T_1114; // @[LZD.scala 49:25]
  wire  _T_1115; // @[LZD.scala 49:47]
  wire  _T_1116; // @[LZD.scala 49:59]
  wire  _T_1117; // @[LZD.scala 49:35]
  wire [2:0] _T_1119; // @[Cat.scala 29:58]
  wire  _T_1120; // @[Shift.scala 12:21]
  wire  _T_1121; // @[Shift.scala 12:21]
  wire  _T_1122; // @[LZD.scala 49:16]
  wire  _T_1123; // @[LZD.scala 49:27]
  wire  _T_1124; // @[LZD.scala 49:25]
  wire [1:0] _T_1125; // @[LZD.scala 49:47]
  wire [1:0] _T_1126; // @[LZD.scala 49:59]
  wire [1:0] _T_1127; // @[LZD.scala 49:35]
  wire [3:0] _T_1129; // @[Cat.scala 29:58]
  wire  _T_1130; // @[Shift.scala 12:21]
  wire  _T_1131; // @[Shift.scala 12:21]
  wire  _T_1132; // @[LZD.scala 49:16]
  wire  _T_1133; // @[LZD.scala 49:27]
  wire  _T_1134; // @[LZD.scala 49:25]
  wire [2:0] _T_1135; // @[LZD.scala 49:47]
  wire [2:0] _T_1136; // @[LZD.scala 49:59]
  wire [2:0] _T_1137; // @[LZD.scala 49:35]
  wire [4:0] _T_1139; // @[Cat.scala 29:58]
  wire [15:0] _T_1140; // @[LZD.scala 44:32]
  wire [7:0] _T_1141; // @[LZD.scala 43:32]
  wire [3:0] _T_1142; // @[LZD.scala 43:32]
  wire [1:0] _T_1143; // @[LZD.scala 43:32]
  wire  _T_1144; // @[LZD.scala 39:14]
  wire  _T_1145; // @[LZD.scala 39:21]
  wire  _T_1146; // @[LZD.scala 39:30]
  wire  _T_1147; // @[LZD.scala 39:27]
  wire  _T_1148; // @[LZD.scala 39:25]
  wire [1:0] _T_1149; // @[Cat.scala 29:58]
  wire [1:0] _T_1150; // @[LZD.scala 44:32]
  wire  _T_1151; // @[LZD.scala 39:14]
  wire  _T_1152; // @[LZD.scala 39:21]
  wire  _T_1153; // @[LZD.scala 39:30]
  wire  _T_1154; // @[LZD.scala 39:27]
  wire  _T_1155; // @[LZD.scala 39:25]
  wire [1:0] _T_1156; // @[Cat.scala 29:58]
  wire  _T_1157; // @[Shift.scala 12:21]
  wire  _T_1158; // @[Shift.scala 12:21]
  wire  _T_1159; // @[LZD.scala 49:16]
  wire  _T_1160; // @[LZD.scala 49:27]
  wire  _T_1161; // @[LZD.scala 49:25]
  wire  _T_1162; // @[LZD.scala 49:47]
  wire  _T_1163; // @[LZD.scala 49:59]
  wire  _T_1164; // @[LZD.scala 49:35]
  wire [2:0] _T_1166; // @[Cat.scala 29:58]
  wire [3:0] _T_1167; // @[LZD.scala 44:32]
  wire [1:0] _T_1168; // @[LZD.scala 43:32]
  wire  _T_1169; // @[LZD.scala 39:14]
  wire  _T_1170; // @[LZD.scala 39:21]
  wire  _T_1171; // @[LZD.scala 39:30]
  wire  _T_1172; // @[LZD.scala 39:27]
  wire  _T_1173; // @[LZD.scala 39:25]
  wire [1:0] _T_1174; // @[Cat.scala 29:58]
  wire [1:0] _T_1175; // @[LZD.scala 44:32]
  wire  _T_1176; // @[LZD.scala 39:14]
  wire  _T_1177; // @[LZD.scala 39:21]
  wire  _T_1178; // @[LZD.scala 39:30]
  wire  _T_1179; // @[LZD.scala 39:27]
  wire  _T_1180; // @[LZD.scala 39:25]
  wire [1:0] _T_1181; // @[Cat.scala 29:58]
  wire  _T_1182; // @[Shift.scala 12:21]
  wire  _T_1183; // @[Shift.scala 12:21]
  wire  _T_1184; // @[LZD.scala 49:16]
  wire  _T_1185; // @[LZD.scala 49:27]
  wire  _T_1186; // @[LZD.scala 49:25]
  wire  _T_1187; // @[LZD.scala 49:47]
  wire  _T_1188; // @[LZD.scala 49:59]
  wire  _T_1189; // @[LZD.scala 49:35]
  wire [2:0] _T_1191; // @[Cat.scala 29:58]
  wire  _T_1192; // @[Shift.scala 12:21]
  wire  _T_1193; // @[Shift.scala 12:21]
  wire  _T_1194; // @[LZD.scala 49:16]
  wire  _T_1195; // @[LZD.scala 49:27]
  wire  _T_1196; // @[LZD.scala 49:25]
  wire [1:0] _T_1197; // @[LZD.scala 49:47]
  wire [1:0] _T_1198; // @[LZD.scala 49:59]
  wire [1:0] _T_1199; // @[LZD.scala 49:35]
  wire [3:0] _T_1201; // @[Cat.scala 29:58]
  wire [7:0] _T_1202; // @[LZD.scala 44:32]
  wire [3:0] _T_1203; // @[LZD.scala 43:32]
  wire [1:0] _T_1204; // @[LZD.scala 43:32]
  wire  _T_1205; // @[LZD.scala 39:14]
  wire  _T_1206; // @[LZD.scala 39:21]
  wire  _T_1207; // @[LZD.scala 39:30]
  wire  _T_1208; // @[LZD.scala 39:27]
  wire  _T_1209; // @[LZD.scala 39:25]
  wire [1:0] _T_1210; // @[Cat.scala 29:58]
  wire [1:0] _T_1211; // @[LZD.scala 44:32]
  wire  _T_1212; // @[LZD.scala 39:14]
  wire  _T_1213; // @[LZD.scala 39:21]
  wire  _T_1214; // @[LZD.scala 39:30]
  wire  _T_1215; // @[LZD.scala 39:27]
  wire  _T_1216; // @[LZD.scala 39:25]
  wire [1:0] _T_1217; // @[Cat.scala 29:58]
  wire  _T_1218; // @[Shift.scala 12:21]
  wire  _T_1219; // @[Shift.scala 12:21]
  wire  _T_1220; // @[LZD.scala 49:16]
  wire  _T_1221; // @[LZD.scala 49:27]
  wire  _T_1222; // @[LZD.scala 49:25]
  wire  _T_1223; // @[LZD.scala 49:47]
  wire  _T_1224; // @[LZD.scala 49:59]
  wire  _T_1225; // @[LZD.scala 49:35]
  wire [2:0] _T_1227; // @[Cat.scala 29:58]
  wire [3:0] _T_1228; // @[LZD.scala 44:32]
  wire [1:0] _T_1229; // @[LZD.scala 43:32]
  wire  _T_1230; // @[LZD.scala 39:14]
  wire  _T_1231; // @[LZD.scala 39:21]
  wire  _T_1232; // @[LZD.scala 39:30]
  wire  _T_1233; // @[LZD.scala 39:27]
  wire  _T_1234; // @[LZD.scala 39:25]
  wire [1:0] _T_1235; // @[Cat.scala 29:58]
  wire [1:0] _T_1236; // @[LZD.scala 44:32]
  wire  _T_1237; // @[LZD.scala 39:14]
  wire  _T_1238; // @[LZD.scala 39:21]
  wire  _T_1239; // @[LZD.scala 39:30]
  wire  _T_1240; // @[LZD.scala 39:27]
  wire  _T_1241; // @[LZD.scala 39:25]
  wire [1:0] _T_1242; // @[Cat.scala 29:58]
  wire  _T_1243; // @[Shift.scala 12:21]
  wire  _T_1244; // @[Shift.scala 12:21]
  wire  _T_1245; // @[LZD.scala 49:16]
  wire  _T_1246; // @[LZD.scala 49:27]
  wire  _T_1247; // @[LZD.scala 49:25]
  wire  _T_1248; // @[LZD.scala 49:47]
  wire  _T_1249; // @[LZD.scala 49:59]
  wire  _T_1250; // @[LZD.scala 49:35]
  wire [2:0] _T_1252; // @[Cat.scala 29:58]
  wire  _T_1253; // @[Shift.scala 12:21]
  wire  _T_1254; // @[Shift.scala 12:21]
  wire  _T_1255; // @[LZD.scala 49:16]
  wire  _T_1256; // @[LZD.scala 49:27]
  wire  _T_1257; // @[LZD.scala 49:25]
  wire [1:0] _T_1258; // @[LZD.scala 49:47]
  wire [1:0] _T_1259; // @[LZD.scala 49:59]
  wire [1:0] _T_1260; // @[LZD.scala 49:35]
  wire [3:0] _T_1262; // @[Cat.scala 29:58]
  wire  _T_1263; // @[Shift.scala 12:21]
  wire  _T_1264; // @[Shift.scala 12:21]
  wire  _T_1265; // @[LZD.scala 49:16]
  wire  _T_1266; // @[LZD.scala 49:27]
  wire  _T_1267; // @[LZD.scala 49:25]
  wire [2:0] _T_1268; // @[LZD.scala 49:47]
  wire [2:0] _T_1269; // @[LZD.scala 49:59]
  wire [2:0] _T_1270; // @[LZD.scala 49:35]
  wire [4:0] _T_1272; // @[Cat.scala 29:58]
  wire  _T_1273; // @[Shift.scala 12:21]
  wire  _T_1274; // @[Shift.scala 12:21]
  wire  _T_1275; // @[LZD.scala 49:16]
  wire  _T_1276; // @[LZD.scala 49:27]
  wire  _T_1277; // @[LZD.scala 49:25]
  wire [3:0] _T_1278; // @[LZD.scala 49:47]
  wire [3:0] _T_1279; // @[LZD.scala 49:59]
  wire [3:0] _T_1280; // @[LZD.scala 49:35]
  wire [5:0] _T_1282; // @[Cat.scala 29:58]
  wire [16:0] _T_1283; // @[LZD.scala 44:32]
  wire [15:0] _T_1284; // @[LZD.scala 43:32]
  wire [7:0] _T_1285; // @[LZD.scala 43:32]
  wire [3:0] _T_1286; // @[LZD.scala 43:32]
  wire [1:0] _T_1287; // @[LZD.scala 43:32]
  wire  _T_1288; // @[LZD.scala 39:14]
  wire  _T_1289; // @[LZD.scala 39:21]
  wire  _T_1290; // @[LZD.scala 39:30]
  wire  _T_1291; // @[LZD.scala 39:27]
  wire  _T_1292; // @[LZD.scala 39:25]
  wire [1:0] _T_1293; // @[Cat.scala 29:58]
  wire [1:0] _T_1294; // @[LZD.scala 44:32]
  wire  _T_1295; // @[LZD.scala 39:14]
  wire  _T_1296; // @[LZD.scala 39:21]
  wire  _T_1297; // @[LZD.scala 39:30]
  wire  _T_1298; // @[LZD.scala 39:27]
  wire  _T_1299; // @[LZD.scala 39:25]
  wire [1:0] _T_1300; // @[Cat.scala 29:58]
  wire  _T_1301; // @[Shift.scala 12:21]
  wire  _T_1302; // @[Shift.scala 12:21]
  wire  _T_1303; // @[LZD.scala 49:16]
  wire  _T_1304; // @[LZD.scala 49:27]
  wire  _T_1305; // @[LZD.scala 49:25]
  wire  _T_1306; // @[LZD.scala 49:47]
  wire  _T_1307; // @[LZD.scala 49:59]
  wire  _T_1308; // @[LZD.scala 49:35]
  wire [2:0] _T_1310; // @[Cat.scala 29:58]
  wire [3:0] _T_1311; // @[LZD.scala 44:32]
  wire [1:0] _T_1312; // @[LZD.scala 43:32]
  wire  _T_1313; // @[LZD.scala 39:14]
  wire  _T_1314; // @[LZD.scala 39:21]
  wire  _T_1315; // @[LZD.scala 39:30]
  wire  _T_1316; // @[LZD.scala 39:27]
  wire  _T_1317; // @[LZD.scala 39:25]
  wire [1:0] _T_1318; // @[Cat.scala 29:58]
  wire [1:0] _T_1319; // @[LZD.scala 44:32]
  wire  _T_1320; // @[LZD.scala 39:14]
  wire  _T_1321; // @[LZD.scala 39:21]
  wire  _T_1322; // @[LZD.scala 39:30]
  wire  _T_1323; // @[LZD.scala 39:27]
  wire  _T_1324; // @[LZD.scala 39:25]
  wire [1:0] _T_1325; // @[Cat.scala 29:58]
  wire  _T_1326; // @[Shift.scala 12:21]
  wire  _T_1327; // @[Shift.scala 12:21]
  wire  _T_1328; // @[LZD.scala 49:16]
  wire  _T_1329; // @[LZD.scala 49:27]
  wire  _T_1330; // @[LZD.scala 49:25]
  wire  _T_1331; // @[LZD.scala 49:47]
  wire  _T_1332; // @[LZD.scala 49:59]
  wire  _T_1333; // @[LZD.scala 49:35]
  wire [2:0] _T_1335; // @[Cat.scala 29:58]
  wire  _T_1336; // @[Shift.scala 12:21]
  wire  _T_1337; // @[Shift.scala 12:21]
  wire  _T_1338; // @[LZD.scala 49:16]
  wire  _T_1339; // @[LZD.scala 49:27]
  wire  _T_1340; // @[LZD.scala 49:25]
  wire [1:0] _T_1341; // @[LZD.scala 49:47]
  wire [1:0] _T_1342; // @[LZD.scala 49:59]
  wire [1:0] _T_1343; // @[LZD.scala 49:35]
  wire [3:0] _T_1345; // @[Cat.scala 29:58]
  wire [7:0] _T_1346; // @[LZD.scala 44:32]
  wire [3:0] _T_1347; // @[LZD.scala 43:32]
  wire [1:0] _T_1348; // @[LZD.scala 43:32]
  wire  _T_1349; // @[LZD.scala 39:14]
  wire  _T_1350; // @[LZD.scala 39:21]
  wire  _T_1351; // @[LZD.scala 39:30]
  wire  _T_1352; // @[LZD.scala 39:27]
  wire  _T_1353; // @[LZD.scala 39:25]
  wire [1:0] _T_1354; // @[Cat.scala 29:58]
  wire [1:0] _T_1355; // @[LZD.scala 44:32]
  wire  _T_1356; // @[LZD.scala 39:14]
  wire  _T_1357; // @[LZD.scala 39:21]
  wire  _T_1358; // @[LZD.scala 39:30]
  wire  _T_1359; // @[LZD.scala 39:27]
  wire  _T_1360; // @[LZD.scala 39:25]
  wire [1:0] _T_1361; // @[Cat.scala 29:58]
  wire  _T_1362; // @[Shift.scala 12:21]
  wire  _T_1363; // @[Shift.scala 12:21]
  wire  _T_1364; // @[LZD.scala 49:16]
  wire  _T_1365; // @[LZD.scala 49:27]
  wire  _T_1366; // @[LZD.scala 49:25]
  wire  _T_1367; // @[LZD.scala 49:47]
  wire  _T_1368; // @[LZD.scala 49:59]
  wire  _T_1369; // @[LZD.scala 49:35]
  wire [2:0] _T_1371; // @[Cat.scala 29:58]
  wire [3:0] _T_1372; // @[LZD.scala 44:32]
  wire [1:0] _T_1373; // @[LZD.scala 43:32]
  wire  _T_1374; // @[LZD.scala 39:14]
  wire  _T_1375; // @[LZD.scala 39:21]
  wire  _T_1376; // @[LZD.scala 39:30]
  wire  _T_1377; // @[LZD.scala 39:27]
  wire  _T_1378; // @[LZD.scala 39:25]
  wire [1:0] _T_1379; // @[Cat.scala 29:58]
  wire [1:0] _T_1380; // @[LZD.scala 44:32]
  wire  _T_1381; // @[LZD.scala 39:14]
  wire  _T_1382; // @[LZD.scala 39:21]
  wire  _T_1383; // @[LZD.scala 39:30]
  wire  _T_1384; // @[LZD.scala 39:27]
  wire  _T_1385; // @[LZD.scala 39:25]
  wire [1:0] _T_1386; // @[Cat.scala 29:58]
  wire  _T_1387; // @[Shift.scala 12:21]
  wire  _T_1388; // @[Shift.scala 12:21]
  wire  _T_1389; // @[LZD.scala 49:16]
  wire  _T_1390; // @[LZD.scala 49:27]
  wire  _T_1391; // @[LZD.scala 49:25]
  wire  _T_1392; // @[LZD.scala 49:47]
  wire  _T_1393; // @[LZD.scala 49:59]
  wire  _T_1394; // @[LZD.scala 49:35]
  wire [2:0] _T_1396; // @[Cat.scala 29:58]
  wire  _T_1397; // @[Shift.scala 12:21]
  wire  _T_1398; // @[Shift.scala 12:21]
  wire  _T_1399; // @[LZD.scala 49:16]
  wire  _T_1400; // @[LZD.scala 49:27]
  wire  _T_1401; // @[LZD.scala 49:25]
  wire [1:0] _T_1402; // @[LZD.scala 49:47]
  wire [1:0] _T_1403; // @[LZD.scala 49:59]
  wire [1:0] _T_1404; // @[LZD.scala 49:35]
  wire [3:0] _T_1406; // @[Cat.scala 29:58]
  wire  _T_1407; // @[Shift.scala 12:21]
  wire  _T_1408; // @[Shift.scala 12:21]
  wire  _T_1409; // @[LZD.scala 49:16]
  wire  _T_1410; // @[LZD.scala 49:27]
  wire  _T_1411; // @[LZD.scala 49:25]
  wire [2:0] _T_1412; // @[LZD.scala 49:47]
  wire [2:0] _T_1413; // @[LZD.scala 49:59]
  wire [2:0] _T_1414; // @[LZD.scala 49:35]
  wire [4:0] _T_1416; // @[Cat.scala 29:58]
  wire  _T_1417; // @[LZD.scala 44:32]
  wire  _T_1419; // @[Shift.scala 12:21]
  wire [3:0] _T_1422; // @[Cat.scala 29:58]
  wire [3:0] _T_1423; // @[LZD.scala 55:32]
  wire [3:0] _T_1424; // @[LZD.scala 55:20]
  wire [4:0] _T_1425; // @[Cat.scala 29:58]
  wire  _T_1426; // @[Shift.scala 12:21]
  wire [4:0] _T_1428; // @[LZD.scala 55:32]
  wire [4:0] _T_1429; // @[LZD.scala 55:20]
  wire [5:0] sumLZD; // @[Cat.scala 29:58]
  wire [5:0] shiftValue; // @[PositFMA.scala 127:24]
  wire [47:0] _T_1430; // @[PositFMA.scala 128:38]
  wire  _T_1431; // @[Shift.scala 16:24]
  wire  _T_1433; // @[Shift.scala 12:21]
  wire [15:0] _T_1434; // @[Shift.scala 64:52]
  wire [47:0] _T_1436; // @[Cat.scala 29:58]
  wire [47:0] _T_1437; // @[Shift.scala 64:27]
  wire [4:0] _T_1438; // @[Shift.scala 66:70]
  wire  _T_1439; // @[Shift.scala 12:21]
  wire [31:0] _T_1440; // @[Shift.scala 64:52]
  wire [47:0] _T_1442; // @[Cat.scala 29:58]
  wire [47:0] _T_1443; // @[Shift.scala 64:27]
  wire [3:0] _T_1444; // @[Shift.scala 66:70]
  wire  _T_1445; // @[Shift.scala 12:21]
  wire [39:0] _T_1446; // @[Shift.scala 64:52]
  wire [47:0] _T_1448; // @[Cat.scala 29:58]
  wire [47:0] _T_1449; // @[Shift.scala 64:27]
  wire [2:0] _T_1450; // @[Shift.scala 66:70]
  wire  _T_1451; // @[Shift.scala 12:21]
  wire [43:0] _T_1452; // @[Shift.scala 64:52]
  wire [47:0] _T_1454; // @[Cat.scala 29:58]
  wire [47:0] _T_1455; // @[Shift.scala 64:27]
  wire [1:0] _T_1456; // @[Shift.scala 66:70]
  wire  _T_1457; // @[Shift.scala 12:21]
  wire [45:0] _T_1458; // @[Shift.scala 64:52]
  wire [47:0] _T_1460; // @[Cat.scala 29:58]
  wire [47:0] _T_1461; // @[Shift.scala 64:27]
  wire  _T_1462; // @[Shift.scala 66:70]
  wire [46:0] _T_1464; // @[Shift.scala 64:52]
  wire [47:0] _T_1465; // @[Cat.scala 29:58]
  wire [47:0] _T_1466; // @[Shift.scala 64:27]
  wire [47:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [9:0] _T_1468; // @[PositFMA.scala 131:36]
  wire [9:0] _T_1469; // @[PositFMA.scala 131:36]
  wire [6:0] _T_1470; // @[Cat.scala 29:58]
  wire [6:0] _T_1471; // @[PositFMA.scala 131:61]
  wire [9:0] _GEN_20; // @[PositFMA.scala 131:42]
  wire [9:0] _T_1473; // @[PositFMA.scala 131:42]
  wire [9:0] sumScale; // @[PositFMA.scala 131:42]
  wire [22:0] sumFrac; // @[PositFMA.scala 132:41]
  wire [24:0] grsTmp; // @[PositFMA.scala 135:41]
  wire [1:0] _T_1474; // @[PositFMA.scala 138:40]
  wire [22:0] _T_1475; // @[PositFMA.scala 138:56]
  wire  _T_1476; // @[PositFMA.scala 138:60]
  wire  underflow; // @[PositFMA.scala 145:32]
  wire  overflow; // @[PositFMA.scala 146:32]
  wire  _T_1477; // @[PositFMA.scala 155:32]
  wire  decF_isZero; // @[PositFMA.scala 155:20]
  wire [9:0] _T_1479; // @[Mux.scala 87:16]
  wire [9:0] _T_1480; // @[Mux.scala 87:16]
  wire [8:0] _GEN_21; // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  wire [8:0] decF_scale; // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  wire [2:0] _T_1481; // @[convert.scala 46:61]
  wire [2:0] _T_1482; // @[convert.scala 46:52]
  wire [2:0] _T_1484; // @[convert.scala 46:42]
  wire [5:0] _T_1485; // @[convert.scala 48:34]
  wire  _T_1486; // @[convert.scala 49:36]
  wire [5:0] _T_1488; // @[convert.scala 50:36]
  wire [5:0] _T_1489; // @[convert.scala 50:36]
  wire [5:0] _T_1490; // @[convert.scala 50:28]
  wire  _T_1491; // @[convert.scala 51:31]
  wire  _T_1492; // @[convert.scala 52:43]
  wire [30:0] _T_1496; // @[Cat.scala 29:58]
  wire [5:0] _T_1497; // @[Shift.scala 39:17]
  wire  _T_1498; // @[Shift.scala 39:24]
  wire [4:0] _T_1499; // @[Shift.scala 40:44]
  wire [14:0] _T_1500; // @[Shift.scala 90:30]
  wire [15:0] _T_1501; // @[Shift.scala 90:48]
  wire  _T_1502; // @[Shift.scala 90:57]
  wire [14:0] _GEN_22; // @[Shift.scala 90:39]
  wire [14:0] _T_1503; // @[Shift.scala 90:39]
  wire  _T_1504; // @[Shift.scala 12:21]
  wire  _T_1505; // @[Shift.scala 12:21]
  wire [15:0] _T_1507; // @[Bitwise.scala 71:12]
  wire [30:0] _T_1508; // @[Cat.scala 29:58]
  wire [30:0] _T_1509; // @[Shift.scala 91:22]
  wire [3:0] _T_1510; // @[Shift.scala 92:77]
  wire [22:0] _T_1511; // @[Shift.scala 90:30]
  wire [7:0] _T_1512; // @[Shift.scala 90:48]
  wire  _T_1513; // @[Shift.scala 90:57]
  wire [22:0] _GEN_23; // @[Shift.scala 90:39]
  wire [22:0] _T_1514; // @[Shift.scala 90:39]
  wire  _T_1515; // @[Shift.scala 12:21]
  wire  _T_1516; // @[Shift.scala 12:21]
  wire [7:0] _T_1518; // @[Bitwise.scala 71:12]
  wire [30:0] _T_1519; // @[Cat.scala 29:58]
  wire [30:0] _T_1520; // @[Shift.scala 91:22]
  wire [2:0] _T_1521; // @[Shift.scala 92:77]
  wire [26:0] _T_1522; // @[Shift.scala 90:30]
  wire [3:0] _T_1523; // @[Shift.scala 90:48]
  wire  _T_1524; // @[Shift.scala 90:57]
  wire [26:0] _GEN_24; // @[Shift.scala 90:39]
  wire [26:0] _T_1525; // @[Shift.scala 90:39]
  wire  _T_1526; // @[Shift.scala 12:21]
  wire  _T_1527; // @[Shift.scala 12:21]
  wire [3:0] _T_1529; // @[Bitwise.scala 71:12]
  wire [30:0] _T_1530; // @[Cat.scala 29:58]
  wire [30:0] _T_1531; // @[Shift.scala 91:22]
  wire [1:0] _T_1532; // @[Shift.scala 92:77]
  wire [28:0] _T_1533; // @[Shift.scala 90:30]
  wire [1:0] _T_1534; // @[Shift.scala 90:48]
  wire  _T_1535; // @[Shift.scala 90:57]
  wire [28:0] _GEN_25; // @[Shift.scala 90:39]
  wire [28:0] _T_1536; // @[Shift.scala 90:39]
  wire  _T_1537; // @[Shift.scala 12:21]
  wire  _T_1538; // @[Shift.scala 12:21]
  wire [1:0] _T_1540; // @[Bitwise.scala 71:12]
  wire [30:0] _T_1541; // @[Cat.scala 29:58]
  wire [30:0] _T_1542; // @[Shift.scala 91:22]
  wire  _T_1543; // @[Shift.scala 92:77]
  wire [29:0] _T_1544; // @[Shift.scala 90:30]
  wire  _T_1545; // @[Shift.scala 90:48]
  wire [29:0] _GEN_26; // @[Shift.scala 90:39]
  wire [29:0] _T_1547; // @[Shift.scala 90:39]
  wire  _T_1549; // @[Shift.scala 12:21]
  wire [30:0] _T_1550; // @[Cat.scala 29:58]
  wire [30:0] _T_1551; // @[Shift.scala 91:22]
  wire [30:0] _T_1554; // @[Bitwise.scala 71:12]
  wire [30:0] _T_1555; // @[Shift.scala 39:10]
  wire  _T_1556; // @[convert.scala 55:31]
  wire  _T_1557; // @[convert.scala 56:31]
  wire  _T_1558; // @[convert.scala 57:31]
  wire  _T_1559; // @[convert.scala 58:31]
  wire [27:0] _T_1560; // @[convert.scala 59:69]
  wire  _T_1561; // @[convert.scala 59:81]
  wire  _T_1562; // @[convert.scala 59:50]
  wire  _T_1564; // @[convert.scala 60:81]
  wire  _T_1565; // @[convert.scala 61:44]
  wire  _T_1566; // @[convert.scala 61:52]
  wire  _T_1567; // @[convert.scala 61:36]
  wire  _T_1568; // @[convert.scala 62:63]
  wire  _T_1569; // @[convert.scala 62:103]
  wire  _T_1570; // @[convert.scala 62:60]
  wire [27:0] _GEN_27; // @[convert.scala 63:56]
  wire [27:0] _T_1573; // @[convert.scala 63:56]
  wire [28:0] _T_1574; // @[Cat.scala 29:58]
  reg  _T_1578; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [28:0] _T_1582; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 29'h1fffffff : 29'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{28'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 29'h1fffffff : 29'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{28'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[28]; // @[convert.scala 18:24]
  assign _T_14 = realA[27]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[27:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[26:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[26:11]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[15:8]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20[7:4]; // @[LZD.scala 43:32]
  assign _T_22 = _T_21[3:2]; // @[LZD.scala 43:32]
  assign _T_23 = _T_22 != 2'h0; // @[LZD.scala 39:14]
  assign _T_24 = _T_22[1]; // @[LZD.scala 39:21]
  assign _T_25 = _T_22[0]; // @[LZD.scala 39:30]
  assign _T_26 = ~ _T_25; // @[LZD.scala 39:27]
  assign _T_27 = _T_24 | _T_26; // @[LZD.scala 39:25]
  assign _T_28 = {_T_23,_T_27}; // @[Cat.scala 29:58]
  assign _T_29 = _T_21[1:0]; // @[LZD.scala 44:32]
  assign _T_30 = _T_29 != 2'h0; // @[LZD.scala 39:14]
  assign _T_31 = _T_29[1]; // @[LZD.scala 39:21]
  assign _T_32 = _T_29[0]; // @[LZD.scala 39:30]
  assign _T_33 = ~ _T_32; // @[LZD.scala 39:27]
  assign _T_34 = _T_31 | _T_33; // @[LZD.scala 39:25]
  assign _T_35 = {_T_30,_T_34}; // @[Cat.scala 29:58]
  assign _T_36 = _T_28[1]; // @[Shift.scala 12:21]
  assign _T_37 = _T_35[1]; // @[Shift.scala 12:21]
  assign _T_38 = _T_36 | _T_37; // @[LZD.scala 49:16]
  assign _T_39 = ~ _T_37; // @[LZD.scala 49:27]
  assign _T_40 = _T_36 | _T_39; // @[LZD.scala 49:25]
  assign _T_41 = _T_28[0:0]; // @[LZD.scala 49:47]
  assign _T_42 = _T_35[0:0]; // @[LZD.scala 49:59]
  assign _T_43 = _T_36 ? _T_41 : _T_42; // @[LZD.scala 49:35]
  assign _T_45 = {_T_38,_T_40,_T_43}; // @[Cat.scala 29:58]
  assign _T_46 = _T_20[3:0]; // @[LZD.scala 44:32]
  assign _T_47 = _T_46[3:2]; // @[LZD.scala 43:32]
  assign _T_48 = _T_47 != 2'h0; // @[LZD.scala 39:14]
  assign _T_49 = _T_47[1]; // @[LZD.scala 39:21]
  assign _T_50 = _T_47[0]; // @[LZD.scala 39:30]
  assign _T_51 = ~ _T_50; // @[LZD.scala 39:27]
  assign _T_52 = _T_49 | _T_51; // @[LZD.scala 39:25]
  assign _T_53 = {_T_48,_T_52}; // @[Cat.scala 29:58]
  assign _T_54 = _T_46[1:0]; // @[LZD.scala 44:32]
  assign _T_55 = _T_54 != 2'h0; // @[LZD.scala 39:14]
  assign _T_56 = _T_54[1]; // @[LZD.scala 39:21]
  assign _T_57 = _T_54[0]; // @[LZD.scala 39:30]
  assign _T_58 = ~ _T_57; // @[LZD.scala 39:27]
  assign _T_59 = _T_56 | _T_58; // @[LZD.scala 39:25]
  assign _T_60 = {_T_55,_T_59}; // @[Cat.scala 29:58]
  assign _T_61 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60[1]; // @[Shift.scala 12:21]
  assign _T_63 = _T_61 | _T_62; // @[LZD.scala 49:16]
  assign _T_64 = ~ _T_62; // @[LZD.scala 49:27]
  assign _T_65 = _T_61 | _T_64; // @[LZD.scala 49:25]
  assign _T_66 = _T_53[0:0]; // @[LZD.scala 49:47]
  assign _T_67 = _T_60[0:0]; // @[LZD.scala 49:59]
  assign _T_68 = _T_61 ? _T_66 : _T_67; // @[LZD.scala 49:35]
  assign _T_70 = {_T_63,_T_65,_T_68}; // @[Cat.scala 29:58]
  assign _T_71 = _T_45[2]; // @[Shift.scala 12:21]
  assign _T_72 = _T_70[2]; // @[Shift.scala 12:21]
  assign _T_73 = _T_71 | _T_72; // @[LZD.scala 49:16]
  assign _T_74 = ~ _T_72; // @[LZD.scala 49:27]
  assign _T_75 = _T_71 | _T_74; // @[LZD.scala 49:25]
  assign _T_76 = _T_45[1:0]; // @[LZD.scala 49:47]
  assign _T_77 = _T_70[1:0]; // @[LZD.scala 49:59]
  assign _T_78 = _T_71 ? _T_76 : _T_77; // @[LZD.scala 49:35]
  assign _T_80 = {_T_73,_T_75,_T_78}; // @[Cat.scala 29:58]
  assign _T_81 = _T_19[7:0]; // @[LZD.scala 44:32]
  assign _T_82 = _T_81[7:4]; // @[LZD.scala 43:32]
  assign _T_83 = _T_82[3:2]; // @[LZD.scala 43:32]
  assign _T_84 = _T_83 != 2'h0; // @[LZD.scala 39:14]
  assign _T_85 = _T_83[1]; // @[LZD.scala 39:21]
  assign _T_86 = _T_83[0]; // @[LZD.scala 39:30]
  assign _T_87 = ~ _T_86; // @[LZD.scala 39:27]
  assign _T_88 = _T_85 | _T_87; // @[LZD.scala 39:25]
  assign _T_89 = {_T_84,_T_88}; // @[Cat.scala 29:58]
  assign _T_90 = _T_82[1:0]; // @[LZD.scala 44:32]
  assign _T_91 = _T_90 != 2'h0; // @[LZD.scala 39:14]
  assign _T_92 = _T_90[1]; // @[LZD.scala 39:21]
  assign _T_93 = _T_90[0]; // @[LZD.scala 39:30]
  assign _T_94 = ~ _T_93; // @[LZD.scala 39:27]
  assign _T_95 = _T_92 | _T_94; // @[LZD.scala 39:25]
  assign _T_96 = {_T_91,_T_95}; // @[Cat.scala 29:58]
  assign _T_97 = _T_89[1]; // @[Shift.scala 12:21]
  assign _T_98 = _T_96[1]; // @[Shift.scala 12:21]
  assign _T_99 = _T_97 | _T_98; // @[LZD.scala 49:16]
  assign _T_100 = ~ _T_98; // @[LZD.scala 49:27]
  assign _T_101 = _T_97 | _T_100; // @[LZD.scala 49:25]
  assign _T_102 = _T_89[0:0]; // @[LZD.scala 49:47]
  assign _T_103 = _T_96[0:0]; // @[LZD.scala 49:59]
  assign _T_104 = _T_97 ? _T_102 : _T_103; // @[LZD.scala 49:35]
  assign _T_106 = {_T_99,_T_101,_T_104}; // @[Cat.scala 29:58]
  assign _T_107 = _T_81[3:0]; // @[LZD.scala 44:32]
  assign _T_108 = _T_107[3:2]; // @[LZD.scala 43:32]
  assign _T_109 = _T_108 != 2'h0; // @[LZD.scala 39:14]
  assign _T_110 = _T_108[1]; // @[LZD.scala 39:21]
  assign _T_111 = _T_108[0]; // @[LZD.scala 39:30]
  assign _T_112 = ~ _T_111; // @[LZD.scala 39:27]
  assign _T_113 = _T_110 | _T_112; // @[LZD.scala 39:25]
  assign _T_114 = {_T_109,_T_113}; // @[Cat.scala 29:58]
  assign _T_115 = _T_107[1:0]; // @[LZD.scala 44:32]
  assign _T_116 = _T_115 != 2'h0; // @[LZD.scala 39:14]
  assign _T_117 = _T_115[1]; // @[LZD.scala 39:21]
  assign _T_118 = _T_115[0]; // @[LZD.scala 39:30]
  assign _T_119 = ~ _T_118; // @[LZD.scala 39:27]
  assign _T_120 = _T_117 | _T_119; // @[LZD.scala 39:25]
  assign _T_121 = {_T_116,_T_120}; // @[Cat.scala 29:58]
  assign _T_122 = _T_114[1]; // @[Shift.scala 12:21]
  assign _T_123 = _T_121[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_122 | _T_123; // @[LZD.scala 49:16]
  assign _T_125 = ~ _T_123; // @[LZD.scala 49:27]
  assign _T_126 = _T_122 | _T_125; // @[LZD.scala 49:25]
  assign _T_127 = _T_114[0:0]; // @[LZD.scala 49:47]
  assign _T_128 = _T_121[0:0]; // @[LZD.scala 49:59]
  assign _T_129 = _T_122 ? _T_127 : _T_128; // @[LZD.scala 49:35]
  assign _T_131 = {_T_124,_T_126,_T_129}; // @[Cat.scala 29:58]
  assign _T_132 = _T_106[2]; // @[Shift.scala 12:21]
  assign _T_133 = _T_131[2]; // @[Shift.scala 12:21]
  assign _T_134 = _T_132 | _T_133; // @[LZD.scala 49:16]
  assign _T_135 = ~ _T_133; // @[LZD.scala 49:27]
  assign _T_136 = _T_132 | _T_135; // @[LZD.scala 49:25]
  assign _T_137 = _T_106[1:0]; // @[LZD.scala 49:47]
  assign _T_138 = _T_131[1:0]; // @[LZD.scala 49:59]
  assign _T_139 = _T_132 ? _T_137 : _T_138; // @[LZD.scala 49:35]
  assign _T_141 = {_T_134,_T_136,_T_139}; // @[Cat.scala 29:58]
  assign _T_142 = _T_80[3]; // @[Shift.scala 12:21]
  assign _T_143 = _T_141[3]; // @[Shift.scala 12:21]
  assign _T_144 = _T_142 | _T_143; // @[LZD.scala 49:16]
  assign _T_145 = ~ _T_143; // @[LZD.scala 49:27]
  assign _T_146 = _T_142 | _T_145; // @[LZD.scala 49:25]
  assign _T_147 = _T_80[2:0]; // @[LZD.scala 49:47]
  assign _T_148 = _T_141[2:0]; // @[LZD.scala 49:59]
  assign _T_149 = _T_142 ? _T_147 : _T_148; // @[LZD.scala 49:35]
  assign _T_151 = {_T_144,_T_146,_T_149}; // @[Cat.scala 29:58]
  assign _T_152 = _T_18[10:0]; // @[LZD.scala 44:32]
  assign _T_153 = _T_152[10:3]; // @[LZD.scala 43:32]
  assign _T_154 = _T_153[7:4]; // @[LZD.scala 43:32]
  assign _T_155 = _T_154[3:2]; // @[LZD.scala 43:32]
  assign _T_156 = _T_155 != 2'h0; // @[LZD.scala 39:14]
  assign _T_157 = _T_155[1]; // @[LZD.scala 39:21]
  assign _T_158 = _T_155[0]; // @[LZD.scala 39:30]
  assign _T_159 = ~ _T_158; // @[LZD.scala 39:27]
  assign _T_160 = _T_157 | _T_159; // @[LZD.scala 39:25]
  assign _T_161 = {_T_156,_T_160}; // @[Cat.scala 29:58]
  assign _T_162 = _T_154[1:0]; // @[LZD.scala 44:32]
  assign _T_163 = _T_162 != 2'h0; // @[LZD.scala 39:14]
  assign _T_164 = _T_162[1]; // @[LZD.scala 39:21]
  assign _T_165 = _T_162[0]; // @[LZD.scala 39:30]
  assign _T_166 = ~ _T_165; // @[LZD.scala 39:27]
  assign _T_167 = _T_164 | _T_166; // @[LZD.scala 39:25]
  assign _T_168 = {_T_163,_T_167}; // @[Cat.scala 29:58]
  assign _T_169 = _T_161[1]; // @[Shift.scala 12:21]
  assign _T_170 = _T_168[1]; // @[Shift.scala 12:21]
  assign _T_171 = _T_169 | _T_170; // @[LZD.scala 49:16]
  assign _T_172 = ~ _T_170; // @[LZD.scala 49:27]
  assign _T_173 = _T_169 | _T_172; // @[LZD.scala 49:25]
  assign _T_174 = _T_161[0:0]; // @[LZD.scala 49:47]
  assign _T_175 = _T_168[0:0]; // @[LZD.scala 49:59]
  assign _T_176 = _T_169 ? _T_174 : _T_175; // @[LZD.scala 49:35]
  assign _T_178 = {_T_171,_T_173,_T_176}; // @[Cat.scala 29:58]
  assign _T_179 = _T_153[3:0]; // @[LZD.scala 44:32]
  assign _T_180 = _T_179[3:2]; // @[LZD.scala 43:32]
  assign _T_181 = _T_180 != 2'h0; // @[LZD.scala 39:14]
  assign _T_182 = _T_180[1]; // @[LZD.scala 39:21]
  assign _T_183 = _T_180[0]; // @[LZD.scala 39:30]
  assign _T_184 = ~ _T_183; // @[LZD.scala 39:27]
  assign _T_185 = _T_182 | _T_184; // @[LZD.scala 39:25]
  assign _T_186 = {_T_181,_T_185}; // @[Cat.scala 29:58]
  assign _T_187 = _T_179[1:0]; // @[LZD.scala 44:32]
  assign _T_188 = _T_187 != 2'h0; // @[LZD.scala 39:14]
  assign _T_189 = _T_187[1]; // @[LZD.scala 39:21]
  assign _T_190 = _T_187[0]; // @[LZD.scala 39:30]
  assign _T_191 = ~ _T_190; // @[LZD.scala 39:27]
  assign _T_192 = _T_189 | _T_191; // @[LZD.scala 39:25]
  assign _T_193 = {_T_188,_T_192}; // @[Cat.scala 29:58]
  assign _T_194 = _T_186[1]; // @[Shift.scala 12:21]
  assign _T_195 = _T_193[1]; // @[Shift.scala 12:21]
  assign _T_196 = _T_194 | _T_195; // @[LZD.scala 49:16]
  assign _T_197 = ~ _T_195; // @[LZD.scala 49:27]
  assign _T_198 = _T_194 | _T_197; // @[LZD.scala 49:25]
  assign _T_199 = _T_186[0:0]; // @[LZD.scala 49:47]
  assign _T_200 = _T_193[0:0]; // @[LZD.scala 49:59]
  assign _T_201 = _T_194 ? _T_199 : _T_200; // @[LZD.scala 49:35]
  assign _T_203 = {_T_196,_T_198,_T_201}; // @[Cat.scala 29:58]
  assign _T_204 = _T_178[2]; // @[Shift.scala 12:21]
  assign _T_205 = _T_203[2]; // @[Shift.scala 12:21]
  assign _T_206 = _T_204 | _T_205; // @[LZD.scala 49:16]
  assign _T_207 = ~ _T_205; // @[LZD.scala 49:27]
  assign _T_208 = _T_204 | _T_207; // @[LZD.scala 49:25]
  assign _T_209 = _T_178[1:0]; // @[LZD.scala 49:47]
  assign _T_210 = _T_203[1:0]; // @[LZD.scala 49:59]
  assign _T_211 = _T_204 ? _T_209 : _T_210; // @[LZD.scala 49:35]
  assign _T_213 = {_T_206,_T_208,_T_211}; // @[Cat.scala 29:58]
  assign _T_214 = _T_152[2:0]; // @[LZD.scala 44:32]
  assign _T_215 = _T_214[2:1]; // @[LZD.scala 43:32]
  assign _T_216 = _T_215 != 2'h0; // @[LZD.scala 39:14]
  assign _T_217 = _T_215[1]; // @[LZD.scala 39:21]
  assign _T_218 = _T_215[0]; // @[LZD.scala 39:30]
  assign _T_219 = ~ _T_218; // @[LZD.scala 39:27]
  assign _T_220 = _T_217 | _T_219; // @[LZD.scala 39:25]
  assign _T_221 = {_T_216,_T_220}; // @[Cat.scala 29:58]
  assign _T_222 = _T_214[0:0]; // @[LZD.scala 44:32]
  assign _T_224 = _T_221[1]; // @[Shift.scala 12:21]
  assign _T_226 = _T_221[0:0]; // @[LZD.scala 55:32]
  assign _T_227 = _T_224 ? _T_226 : _T_222; // @[LZD.scala 55:20]
  assign _T_229 = _T_213[3]; // @[Shift.scala 12:21]
  assign _T_231 = {1'h1,_T_224,_T_227}; // @[Cat.scala 29:58]
  assign _T_232 = _T_213[2:0]; // @[LZD.scala 55:32]
  assign _T_233 = _T_229 ? _T_232 : _T_231; // @[LZD.scala 55:20]
  assign _T_234 = {_T_229,_T_233}; // @[Cat.scala 29:58]
  assign _T_235 = _T_151[4]; // @[Shift.scala 12:21]
  assign _T_237 = _T_151[3:0]; // @[LZD.scala 55:32]
  assign _T_238 = _T_235 ? _T_237 : _T_234; // @[LZD.scala 55:20]
  assign _T_239 = {_T_235,_T_238}; // @[Cat.scala 29:58]
  assign _T_240 = ~ _T_239; // @[convert.scala 21:22]
  assign _T_241 = realA[25:0]; // @[convert.scala 22:36]
  assign _T_242 = _T_240 < 5'h1a; // @[Shift.scala 16:24]
  assign _T_244 = _T_240[4]; // @[Shift.scala 12:21]
  assign _T_245 = _T_241[9:0]; // @[Shift.scala 64:52]
  assign _T_247 = {_T_245,16'h0}; // @[Cat.scala 29:58]
  assign _T_248 = _T_244 ? _T_247 : _T_241; // @[Shift.scala 64:27]
  assign _T_249 = _T_240[3:0]; // @[Shift.scala 66:70]
  assign _T_250 = _T_249[3]; // @[Shift.scala 12:21]
  assign _T_251 = _T_248[17:0]; // @[Shift.scala 64:52]
  assign _T_253 = {_T_251,8'h0}; // @[Cat.scala 29:58]
  assign _T_254 = _T_250 ? _T_253 : _T_248; // @[Shift.scala 64:27]
  assign _T_255 = _T_249[2:0]; // @[Shift.scala 66:70]
  assign _T_256 = _T_255[2]; // @[Shift.scala 12:21]
  assign _T_257 = _T_254[21:0]; // @[Shift.scala 64:52]
  assign _T_259 = {_T_257,4'h0}; // @[Cat.scala 29:58]
  assign _T_260 = _T_256 ? _T_259 : _T_254; // @[Shift.scala 64:27]
  assign _T_261 = _T_255[1:0]; // @[Shift.scala 66:70]
  assign _T_262 = _T_261[1]; // @[Shift.scala 12:21]
  assign _T_263 = _T_260[23:0]; // @[Shift.scala 64:52]
  assign _T_265 = {_T_263,2'h0}; // @[Cat.scala 29:58]
  assign _T_266 = _T_262 ? _T_265 : _T_260; // @[Shift.scala 64:27]
  assign _T_267 = _T_261[0:0]; // @[Shift.scala 66:70]
  assign _T_269 = _T_266[24:0]; // @[Shift.scala 64:52]
  assign _T_270 = {_T_269,1'h0}; // @[Cat.scala 29:58]
  assign _T_271 = _T_267 ? _T_270 : _T_266; // @[Shift.scala 64:27]
  assign _T_272 = _T_242 ? _T_271 : 26'h0; // @[Shift.scala 16:10]
  assign _T_273 = _T_272[25:23]; // @[convert.scala 23:34]
  assign decA_fraction = _T_272[22:0]; // @[convert.scala 24:34]
  assign _T_275 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_277 = _T_15 ? _T_240 : _T_239; // @[convert.scala 25:42]
  assign _T_280 = ~ _T_273; // @[convert.scala 26:67]
  assign _T_281 = _T_13 ? _T_280 : _T_273; // @[convert.scala 26:51]
  assign _T_282 = {_T_275,_T_277,_T_281}; // @[Cat.scala 29:58]
  assign _T_284 = realA[27:0]; // @[convert.scala 29:56]
  assign _T_285 = _T_284 != 28'h0; // @[convert.scala 29:60]
  assign _T_286 = ~ _T_285; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_286; // @[convert.scala 29:39]
  assign _T_289 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_289 & _T_286; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_282); // @[convert.scala 32:24]
  assign _T_298 = io_B[28]; // @[convert.scala 18:24]
  assign _T_299 = io_B[27]; // @[convert.scala 18:40]
  assign _T_300 = _T_298 ^ _T_299; // @[convert.scala 18:36]
  assign _T_301 = io_B[27:1]; // @[convert.scala 19:24]
  assign _T_302 = io_B[26:0]; // @[convert.scala 19:43]
  assign _T_303 = _T_301 ^ _T_302; // @[convert.scala 19:39]
  assign _T_304 = _T_303[26:11]; // @[LZD.scala 43:32]
  assign _T_305 = _T_304[15:8]; // @[LZD.scala 43:32]
  assign _T_306 = _T_305[7:4]; // @[LZD.scala 43:32]
  assign _T_307 = _T_306[3:2]; // @[LZD.scala 43:32]
  assign _T_308 = _T_307 != 2'h0; // @[LZD.scala 39:14]
  assign _T_309 = _T_307[1]; // @[LZD.scala 39:21]
  assign _T_310 = _T_307[0]; // @[LZD.scala 39:30]
  assign _T_311 = ~ _T_310; // @[LZD.scala 39:27]
  assign _T_312 = _T_309 | _T_311; // @[LZD.scala 39:25]
  assign _T_313 = {_T_308,_T_312}; // @[Cat.scala 29:58]
  assign _T_314 = _T_306[1:0]; // @[LZD.scala 44:32]
  assign _T_315 = _T_314 != 2'h0; // @[LZD.scala 39:14]
  assign _T_316 = _T_314[1]; // @[LZD.scala 39:21]
  assign _T_317 = _T_314[0]; // @[LZD.scala 39:30]
  assign _T_318 = ~ _T_317; // @[LZD.scala 39:27]
  assign _T_319 = _T_316 | _T_318; // @[LZD.scala 39:25]
  assign _T_320 = {_T_315,_T_319}; // @[Cat.scala 29:58]
  assign _T_321 = _T_313[1]; // @[Shift.scala 12:21]
  assign _T_322 = _T_320[1]; // @[Shift.scala 12:21]
  assign _T_323 = _T_321 | _T_322; // @[LZD.scala 49:16]
  assign _T_324 = ~ _T_322; // @[LZD.scala 49:27]
  assign _T_325 = _T_321 | _T_324; // @[LZD.scala 49:25]
  assign _T_326 = _T_313[0:0]; // @[LZD.scala 49:47]
  assign _T_327 = _T_320[0:0]; // @[LZD.scala 49:59]
  assign _T_328 = _T_321 ? _T_326 : _T_327; // @[LZD.scala 49:35]
  assign _T_330 = {_T_323,_T_325,_T_328}; // @[Cat.scala 29:58]
  assign _T_331 = _T_305[3:0]; // @[LZD.scala 44:32]
  assign _T_332 = _T_331[3:2]; // @[LZD.scala 43:32]
  assign _T_333 = _T_332 != 2'h0; // @[LZD.scala 39:14]
  assign _T_334 = _T_332[1]; // @[LZD.scala 39:21]
  assign _T_335 = _T_332[0]; // @[LZD.scala 39:30]
  assign _T_336 = ~ _T_335; // @[LZD.scala 39:27]
  assign _T_337 = _T_334 | _T_336; // @[LZD.scala 39:25]
  assign _T_338 = {_T_333,_T_337}; // @[Cat.scala 29:58]
  assign _T_339 = _T_331[1:0]; // @[LZD.scala 44:32]
  assign _T_340 = _T_339 != 2'h0; // @[LZD.scala 39:14]
  assign _T_341 = _T_339[1]; // @[LZD.scala 39:21]
  assign _T_342 = _T_339[0]; // @[LZD.scala 39:30]
  assign _T_343 = ~ _T_342; // @[LZD.scala 39:27]
  assign _T_344 = _T_341 | _T_343; // @[LZD.scala 39:25]
  assign _T_345 = {_T_340,_T_344}; // @[Cat.scala 29:58]
  assign _T_346 = _T_338[1]; // @[Shift.scala 12:21]
  assign _T_347 = _T_345[1]; // @[Shift.scala 12:21]
  assign _T_348 = _T_346 | _T_347; // @[LZD.scala 49:16]
  assign _T_349 = ~ _T_347; // @[LZD.scala 49:27]
  assign _T_350 = _T_346 | _T_349; // @[LZD.scala 49:25]
  assign _T_351 = _T_338[0:0]; // @[LZD.scala 49:47]
  assign _T_352 = _T_345[0:0]; // @[LZD.scala 49:59]
  assign _T_353 = _T_346 ? _T_351 : _T_352; // @[LZD.scala 49:35]
  assign _T_355 = {_T_348,_T_350,_T_353}; // @[Cat.scala 29:58]
  assign _T_356 = _T_330[2]; // @[Shift.scala 12:21]
  assign _T_357 = _T_355[2]; // @[Shift.scala 12:21]
  assign _T_358 = _T_356 | _T_357; // @[LZD.scala 49:16]
  assign _T_359 = ~ _T_357; // @[LZD.scala 49:27]
  assign _T_360 = _T_356 | _T_359; // @[LZD.scala 49:25]
  assign _T_361 = _T_330[1:0]; // @[LZD.scala 49:47]
  assign _T_362 = _T_355[1:0]; // @[LZD.scala 49:59]
  assign _T_363 = _T_356 ? _T_361 : _T_362; // @[LZD.scala 49:35]
  assign _T_365 = {_T_358,_T_360,_T_363}; // @[Cat.scala 29:58]
  assign _T_366 = _T_304[7:0]; // @[LZD.scala 44:32]
  assign _T_367 = _T_366[7:4]; // @[LZD.scala 43:32]
  assign _T_368 = _T_367[3:2]; // @[LZD.scala 43:32]
  assign _T_369 = _T_368 != 2'h0; // @[LZD.scala 39:14]
  assign _T_370 = _T_368[1]; // @[LZD.scala 39:21]
  assign _T_371 = _T_368[0]; // @[LZD.scala 39:30]
  assign _T_372 = ~ _T_371; // @[LZD.scala 39:27]
  assign _T_373 = _T_370 | _T_372; // @[LZD.scala 39:25]
  assign _T_374 = {_T_369,_T_373}; // @[Cat.scala 29:58]
  assign _T_375 = _T_367[1:0]; // @[LZD.scala 44:32]
  assign _T_376 = _T_375 != 2'h0; // @[LZD.scala 39:14]
  assign _T_377 = _T_375[1]; // @[LZD.scala 39:21]
  assign _T_378 = _T_375[0]; // @[LZD.scala 39:30]
  assign _T_379 = ~ _T_378; // @[LZD.scala 39:27]
  assign _T_380 = _T_377 | _T_379; // @[LZD.scala 39:25]
  assign _T_381 = {_T_376,_T_380}; // @[Cat.scala 29:58]
  assign _T_382 = _T_374[1]; // @[Shift.scala 12:21]
  assign _T_383 = _T_381[1]; // @[Shift.scala 12:21]
  assign _T_384 = _T_382 | _T_383; // @[LZD.scala 49:16]
  assign _T_385 = ~ _T_383; // @[LZD.scala 49:27]
  assign _T_386 = _T_382 | _T_385; // @[LZD.scala 49:25]
  assign _T_387 = _T_374[0:0]; // @[LZD.scala 49:47]
  assign _T_388 = _T_381[0:0]; // @[LZD.scala 49:59]
  assign _T_389 = _T_382 ? _T_387 : _T_388; // @[LZD.scala 49:35]
  assign _T_391 = {_T_384,_T_386,_T_389}; // @[Cat.scala 29:58]
  assign _T_392 = _T_366[3:0]; // @[LZD.scala 44:32]
  assign _T_393 = _T_392[3:2]; // @[LZD.scala 43:32]
  assign _T_394 = _T_393 != 2'h0; // @[LZD.scala 39:14]
  assign _T_395 = _T_393[1]; // @[LZD.scala 39:21]
  assign _T_396 = _T_393[0]; // @[LZD.scala 39:30]
  assign _T_397 = ~ _T_396; // @[LZD.scala 39:27]
  assign _T_398 = _T_395 | _T_397; // @[LZD.scala 39:25]
  assign _T_399 = {_T_394,_T_398}; // @[Cat.scala 29:58]
  assign _T_400 = _T_392[1:0]; // @[LZD.scala 44:32]
  assign _T_401 = _T_400 != 2'h0; // @[LZD.scala 39:14]
  assign _T_402 = _T_400[1]; // @[LZD.scala 39:21]
  assign _T_403 = _T_400[0]; // @[LZD.scala 39:30]
  assign _T_404 = ~ _T_403; // @[LZD.scala 39:27]
  assign _T_405 = _T_402 | _T_404; // @[LZD.scala 39:25]
  assign _T_406 = {_T_401,_T_405}; // @[Cat.scala 29:58]
  assign _T_407 = _T_399[1]; // @[Shift.scala 12:21]
  assign _T_408 = _T_406[1]; // @[Shift.scala 12:21]
  assign _T_409 = _T_407 | _T_408; // @[LZD.scala 49:16]
  assign _T_410 = ~ _T_408; // @[LZD.scala 49:27]
  assign _T_411 = _T_407 | _T_410; // @[LZD.scala 49:25]
  assign _T_412 = _T_399[0:0]; // @[LZD.scala 49:47]
  assign _T_413 = _T_406[0:0]; // @[LZD.scala 49:59]
  assign _T_414 = _T_407 ? _T_412 : _T_413; // @[LZD.scala 49:35]
  assign _T_416 = {_T_409,_T_411,_T_414}; // @[Cat.scala 29:58]
  assign _T_417 = _T_391[2]; // @[Shift.scala 12:21]
  assign _T_418 = _T_416[2]; // @[Shift.scala 12:21]
  assign _T_419 = _T_417 | _T_418; // @[LZD.scala 49:16]
  assign _T_420 = ~ _T_418; // @[LZD.scala 49:27]
  assign _T_421 = _T_417 | _T_420; // @[LZD.scala 49:25]
  assign _T_422 = _T_391[1:0]; // @[LZD.scala 49:47]
  assign _T_423 = _T_416[1:0]; // @[LZD.scala 49:59]
  assign _T_424 = _T_417 ? _T_422 : _T_423; // @[LZD.scala 49:35]
  assign _T_426 = {_T_419,_T_421,_T_424}; // @[Cat.scala 29:58]
  assign _T_427 = _T_365[3]; // @[Shift.scala 12:21]
  assign _T_428 = _T_426[3]; // @[Shift.scala 12:21]
  assign _T_429 = _T_427 | _T_428; // @[LZD.scala 49:16]
  assign _T_430 = ~ _T_428; // @[LZD.scala 49:27]
  assign _T_431 = _T_427 | _T_430; // @[LZD.scala 49:25]
  assign _T_432 = _T_365[2:0]; // @[LZD.scala 49:47]
  assign _T_433 = _T_426[2:0]; // @[LZD.scala 49:59]
  assign _T_434 = _T_427 ? _T_432 : _T_433; // @[LZD.scala 49:35]
  assign _T_436 = {_T_429,_T_431,_T_434}; // @[Cat.scala 29:58]
  assign _T_437 = _T_303[10:0]; // @[LZD.scala 44:32]
  assign _T_438 = _T_437[10:3]; // @[LZD.scala 43:32]
  assign _T_439 = _T_438[7:4]; // @[LZD.scala 43:32]
  assign _T_440 = _T_439[3:2]; // @[LZD.scala 43:32]
  assign _T_441 = _T_440 != 2'h0; // @[LZD.scala 39:14]
  assign _T_442 = _T_440[1]; // @[LZD.scala 39:21]
  assign _T_443 = _T_440[0]; // @[LZD.scala 39:30]
  assign _T_444 = ~ _T_443; // @[LZD.scala 39:27]
  assign _T_445 = _T_442 | _T_444; // @[LZD.scala 39:25]
  assign _T_446 = {_T_441,_T_445}; // @[Cat.scala 29:58]
  assign _T_447 = _T_439[1:0]; // @[LZD.scala 44:32]
  assign _T_448 = _T_447 != 2'h0; // @[LZD.scala 39:14]
  assign _T_449 = _T_447[1]; // @[LZD.scala 39:21]
  assign _T_450 = _T_447[0]; // @[LZD.scala 39:30]
  assign _T_451 = ~ _T_450; // @[LZD.scala 39:27]
  assign _T_452 = _T_449 | _T_451; // @[LZD.scala 39:25]
  assign _T_453 = {_T_448,_T_452}; // @[Cat.scala 29:58]
  assign _T_454 = _T_446[1]; // @[Shift.scala 12:21]
  assign _T_455 = _T_453[1]; // @[Shift.scala 12:21]
  assign _T_456 = _T_454 | _T_455; // @[LZD.scala 49:16]
  assign _T_457 = ~ _T_455; // @[LZD.scala 49:27]
  assign _T_458 = _T_454 | _T_457; // @[LZD.scala 49:25]
  assign _T_459 = _T_446[0:0]; // @[LZD.scala 49:47]
  assign _T_460 = _T_453[0:0]; // @[LZD.scala 49:59]
  assign _T_461 = _T_454 ? _T_459 : _T_460; // @[LZD.scala 49:35]
  assign _T_463 = {_T_456,_T_458,_T_461}; // @[Cat.scala 29:58]
  assign _T_464 = _T_438[3:0]; // @[LZD.scala 44:32]
  assign _T_465 = _T_464[3:2]; // @[LZD.scala 43:32]
  assign _T_466 = _T_465 != 2'h0; // @[LZD.scala 39:14]
  assign _T_467 = _T_465[1]; // @[LZD.scala 39:21]
  assign _T_468 = _T_465[0]; // @[LZD.scala 39:30]
  assign _T_469 = ~ _T_468; // @[LZD.scala 39:27]
  assign _T_470 = _T_467 | _T_469; // @[LZD.scala 39:25]
  assign _T_471 = {_T_466,_T_470}; // @[Cat.scala 29:58]
  assign _T_472 = _T_464[1:0]; // @[LZD.scala 44:32]
  assign _T_473 = _T_472 != 2'h0; // @[LZD.scala 39:14]
  assign _T_474 = _T_472[1]; // @[LZD.scala 39:21]
  assign _T_475 = _T_472[0]; // @[LZD.scala 39:30]
  assign _T_476 = ~ _T_475; // @[LZD.scala 39:27]
  assign _T_477 = _T_474 | _T_476; // @[LZD.scala 39:25]
  assign _T_478 = {_T_473,_T_477}; // @[Cat.scala 29:58]
  assign _T_479 = _T_471[1]; // @[Shift.scala 12:21]
  assign _T_480 = _T_478[1]; // @[Shift.scala 12:21]
  assign _T_481 = _T_479 | _T_480; // @[LZD.scala 49:16]
  assign _T_482 = ~ _T_480; // @[LZD.scala 49:27]
  assign _T_483 = _T_479 | _T_482; // @[LZD.scala 49:25]
  assign _T_484 = _T_471[0:0]; // @[LZD.scala 49:47]
  assign _T_485 = _T_478[0:0]; // @[LZD.scala 49:59]
  assign _T_486 = _T_479 ? _T_484 : _T_485; // @[LZD.scala 49:35]
  assign _T_488 = {_T_481,_T_483,_T_486}; // @[Cat.scala 29:58]
  assign _T_489 = _T_463[2]; // @[Shift.scala 12:21]
  assign _T_490 = _T_488[2]; // @[Shift.scala 12:21]
  assign _T_491 = _T_489 | _T_490; // @[LZD.scala 49:16]
  assign _T_492 = ~ _T_490; // @[LZD.scala 49:27]
  assign _T_493 = _T_489 | _T_492; // @[LZD.scala 49:25]
  assign _T_494 = _T_463[1:0]; // @[LZD.scala 49:47]
  assign _T_495 = _T_488[1:0]; // @[LZD.scala 49:59]
  assign _T_496 = _T_489 ? _T_494 : _T_495; // @[LZD.scala 49:35]
  assign _T_498 = {_T_491,_T_493,_T_496}; // @[Cat.scala 29:58]
  assign _T_499 = _T_437[2:0]; // @[LZD.scala 44:32]
  assign _T_500 = _T_499[2:1]; // @[LZD.scala 43:32]
  assign _T_501 = _T_500 != 2'h0; // @[LZD.scala 39:14]
  assign _T_502 = _T_500[1]; // @[LZD.scala 39:21]
  assign _T_503 = _T_500[0]; // @[LZD.scala 39:30]
  assign _T_504 = ~ _T_503; // @[LZD.scala 39:27]
  assign _T_505 = _T_502 | _T_504; // @[LZD.scala 39:25]
  assign _T_506 = {_T_501,_T_505}; // @[Cat.scala 29:58]
  assign _T_507 = _T_499[0:0]; // @[LZD.scala 44:32]
  assign _T_509 = _T_506[1]; // @[Shift.scala 12:21]
  assign _T_511 = _T_506[0:0]; // @[LZD.scala 55:32]
  assign _T_512 = _T_509 ? _T_511 : _T_507; // @[LZD.scala 55:20]
  assign _T_514 = _T_498[3]; // @[Shift.scala 12:21]
  assign _T_516 = {1'h1,_T_509,_T_512}; // @[Cat.scala 29:58]
  assign _T_517 = _T_498[2:0]; // @[LZD.scala 55:32]
  assign _T_518 = _T_514 ? _T_517 : _T_516; // @[LZD.scala 55:20]
  assign _T_519 = {_T_514,_T_518}; // @[Cat.scala 29:58]
  assign _T_520 = _T_436[4]; // @[Shift.scala 12:21]
  assign _T_522 = _T_436[3:0]; // @[LZD.scala 55:32]
  assign _T_523 = _T_520 ? _T_522 : _T_519; // @[LZD.scala 55:20]
  assign _T_524 = {_T_520,_T_523}; // @[Cat.scala 29:58]
  assign _T_525 = ~ _T_524; // @[convert.scala 21:22]
  assign _T_526 = io_B[25:0]; // @[convert.scala 22:36]
  assign _T_527 = _T_525 < 5'h1a; // @[Shift.scala 16:24]
  assign _T_529 = _T_525[4]; // @[Shift.scala 12:21]
  assign _T_530 = _T_526[9:0]; // @[Shift.scala 64:52]
  assign _T_532 = {_T_530,16'h0}; // @[Cat.scala 29:58]
  assign _T_533 = _T_529 ? _T_532 : _T_526; // @[Shift.scala 64:27]
  assign _T_534 = _T_525[3:0]; // @[Shift.scala 66:70]
  assign _T_535 = _T_534[3]; // @[Shift.scala 12:21]
  assign _T_536 = _T_533[17:0]; // @[Shift.scala 64:52]
  assign _T_538 = {_T_536,8'h0}; // @[Cat.scala 29:58]
  assign _T_539 = _T_535 ? _T_538 : _T_533; // @[Shift.scala 64:27]
  assign _T_540 = _T_534[2:0]; // @[Shift.scala 66:70]
  assign _T_541 = _T_540[2]; // @[Shift.scala 12:21]
  assign _T_542 = _T_539[21:0]; // @[Shift.scala 64:52]
  assign _T_544 = {_T_542,4'h0}; // @[Cat.scala 29:58]
  assign _T_545 = _T_541 ? _T_544 : _T_539; // @[Shift.scala 64:27]
  assign _T_546 = _T_540[1:0]; // @[Shift.scala 66:70]
  assign _T_547 = _T_546[1]; // @[Shift.scala 12:21]
  assign _T_548 = _T_545[23:0]; // @[Shift.scala 64:52]
  assign _T_550 = {_T_548,2'h0}; // @[Cat.scala 29:58]
  assign _T_551 = _T_547 ? _T_550 : _T_545; // @[Shift.scala 64:27]
  assign _T_552 = _T_546[0:0]; // @[Shift.scala 66:70]
  assign _T_554 = _T_551[24:0]; // @[Shift.scala 64:52]
  assign _T_555 = {_T_554,1'h0}; // @[Cat.scala 29:58]
  assign _T_556 = _T_552 ? _T_555 : _T_551; // @[Shift.scala 64:27]
  assign _T_557 = _T_527 ? _T_556 : 26'h0; // @[Shift.scala 16:10]
  assign _T_558 = _T_557[25:23]; // @[convert.scala 23:34]
  assign decB_fraction = _T_557[22:0]; // @[convert.scala 24:34]
  assign _T_560 = _T_300 == 1'h0; // @[convert.scala 25:26]
  assign _T_562 = _T_300 ? _T_525 : _T_524; // @[convert.scala 25:42]
  assign _T_565 = ~ _T_558; // @[convert.scala 26:67]
  assign _T_566 = _T_298 ? _T_565 : _T_558; // @[convert.scala 26:51]
  assign _T_567 = {_T_560,_T_562,_T_566}; // @[Cat.scala 29:58]
  assign _T_569 = io_B[27:0]; // @[convert.scala 29:56]
  assign _T_570 = _T_569 != 28'h0; // @[convert.scala 29:60]
  assign _T_571 = ~ _T_570; // @[convert.scala 29:41]
  assign decB_isNaR = _T_298 & _T_571; // @[convert.scala 29:39]
  assign _T_574 = _T_298 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_574 & _T_571; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_567); // @[convert.scala 32:24]
  assign _T_583 = realC[28]; // @[convert.scala 18:24]
  assign _T_584 = realC[27]; // @[convert.scala 18:40]
  assign _T_585 = _T_583 ^ _T_584; // @[convert.scala 18:36]
  assign _T_586 = realC[27:1]; // @[convert.scala 19:24]
  assign _T_587 = realC[26:0]; // @[convert.scala 19:43]
  assign _T_588 = _T_586 ^ _T_587; // @[convert.scala 19:39]
  assign _T_589 = _T_588[26:11]; // @[LZD.scala 43:32]
  assign _T_590 = _T_589[15:8]; // @[LZD.scala 43:32]
  assign _T_591 = _T_590[7:4]; // @[LZD.scala 43:32]
  assign _T_592 = _T_591[3:2]; // @[LZD.scala 43:32]
  assign _T_593 = _T_592 != 2'h0; // @[LZD.scala 39:14]
  assign _T_594 = _T_592[1]; // @[LZD.scala 39:21]
  assign _T_595 = _T_592[0]; // @[LZD.scala 39:30]
  assign _T_596 = ~ _T_595; // @[LZD.scala 39:27]
  assign _T_597 = _T_594 | _T_596; // @[LZD.scala 39:25]
  assign _T_598 = {_T_593,_T_597}; // @[Cat.scala 29:58]
  assign _T_599 = _T_591[1:0]; // @[LZD.scala 44:32]
  assign _T_600 = _T_599 != 2'h0; // @[LZD.scala 39:14]
  assign _T_601 = _T_599[1]; // @[LZD.scala 39:21]
  assign _T_602 = _T_599[0]; // @[LZD.scala 39:30]
  assign _T_603 = ~ _T_602; // @[LZD.scala 39:27]
  assign _T_604 = _T_601 | _T_603; // @[LZD.scala 39:25]
  assign _T_605 = {_T_600,_T_604}; // @[Cat.scala 29:58]
  assign _T_606 = _T_598[1]; // @[Shift.scala 12:21]
  assign _T_607 = _T_605[1]; // @[Shift.scala 12:21]
  assign _T_608 = _T_606 | _T_607; // @[LZD.scala 49:16]
  assign _T_609 = ~ _T_607; // @[LZD.scala 49:27]
  assign _T_610 = _T_606 | _T_609; // @[LZD.scala 49:25]
  assign _T_611 = _T_598[0:0]; // @[LZD.scala 49:47]
  assign _T_612 = _T_605[0:0]; // @[LZD.scala 49:59]
  assign _T_613 = _T_606 ? _T_611 : _T_612; // @[LZD.scala 49:35]
  assign _T_615 = {_T_608,_T_610,_T_613}; // @[Cat.scala 29:58]
  assign _T_616 = _T_590[3:0]; // @[LZD.scala 44:32]
  assign _T_617 = _T_616[3:2]; // @[LZD.scala 43:32]
  assign _T_618 = _T_617 != 2'h0; // @[LZD.scala 39:14]
  assign _T_619 = _T_617[1]; // @[LZD.scala 39:21]
  assign _T_620 = _T_617[0]; // @[LZD.scala 39:30]
  assign _T_621 = ~ _T_620; // @[LZD.scala 39:27]
  assign _T_622 = _T_619 | _T_621; // @[LZD.scala 39:25]
  assign _T_623 = {_T_618,_T_622}; // @[Cat.scala 29:58]
  assign _T_624 = _T_616[1:0]; // @[LZD.scala 44:32]
  assign _T_625 = _T_624 != 2'h0; // @[LZD.scala 39:14]
  assign _T_626 = _T_624[1]; // @[LZD.scala 39:21]
  assign _T_627 = _T_624[0]; // @[LZD.scala 39:30]
  assign _T_628 = ~ _T_627; // @[LZD.scala 39:27]
  assign _T_629 = _T_626 | _T_628; // @[LZD.scala 39:25]
  assign _T_630 = {_T_625,_T_629}; // @[Cat.scala 29:58]
  assign _T_631 = _T_623[1]; // @[Shift.scala 12:21]
  assign _T_632 = _T_630[1]; // @[Shift.scala 12:21]
  assign _T_633 = _T_631 | _T_632; // @[LZD.scala 49:16]
  assign _T_634 = ~ _T_632; // @[LZD.scala 49:27]
  assign _T_635 = _T_631 | _T_634; // @[LZD.scala 49:25]
  assign _T_636 = _T_623[0:0]; // @[LZD.scala 49:47]
  assign _T_637 = _T_630[0:0]; // @[LZD.scala 49:59]
  assign _T_638 = _T_631 ? _T_636 : _T_637; // @[LZD.scala 49:35]
  assign _T_640 = {_T_633,_T_635,_T_638}; // @[Cat.scala 29:58]
  assign _T_641 = _T_615[2]; // @[Shift.scala 12:21]
  assign _T_642 = _T_640[2]; // @[Shift.scala 12:21]
  assign _T_643 = _T_641 | _T_642; // @[LZD.scala 49:16]
  assign _T_644 = ~ _T_642; // @[LZD.scala 49:27]
  assign _T_645 = _T_641 | _T_644; // @[LZD.scala 49:25]
  assign _T_646 = _T_615[1:0]; // @[LZD.scala 49:47]
  assign _T_647 = _T_640[1:0]; // @[LZD.scala 49:59]
  assign _T_648 = _T_641 ? _T_646 : _T_647; // @[LZD.scala 49:35]
  assign _T_650 = {_T_643,_T_645,_T_648}; // @[Cat.scala 29:58]
  assign _T_651 = _T_589[7:0]; // @[LZD.scala 44:32]
  assign _T_652 = _T_651[7:4]; // @[LZD.scala 43:32]
  assign _T_653 = _T_652[3:2]; // @[LZD.scala 43:32]
  assign _T_654 = _T_653 != 2'h0; // @[LZD.scala 39:14]
  assign _T_655 = _T_653[1]; // @[LZD.scala 39:21]
  assign _T_656 = _T_653[0]; // @[LZD.scala 39:30]
  assign _T_657 = ~ _T_656; // @[LZD.scala 39:27]
  assign _T_658 = _T_655 | _T_657; // @[LZD.scala 39:25]
  assign _T_659 = {_T_654,_T_658}; // @[Cat.scala 29:58]
  assign _T_660 = _T_652[1:0]; // @[LZD.scala 44:32]
  assign _T_661 = _T_660 != 2'h0; // @[LZD.scala 39:14]
  assign _T_662 = _T_660[1]; // @[LZD.scala 39:21]
  assign _T_663 = _T_660[0]; // @[LZD.scala 39:30]
  assign _T_664 = ~ _T_663; // @[LZD.scala 39:27]
  assign _T_665 = _T_662 | _T_664; // @[LZD.scala 39:25]
  assign _T_666 = {_T_661,_T_665}; // @[Cat.scala 29:58]
  assign _T_667 = _T_659[1]; // @[Shift.scala 12:21]
  assign _T_668 = _T_666[1]; // @[Shift.scala 12:21]
  assign _T_669 = _T_667 | _T_668; // @[LZD.scala 49:16]
  assign _T_670 = ~ _T_668; // @[LZD.scala 49:27]
  assign _T_671 = _T_667 | _T_670; // @[LZD.scala 49:25]
  assign _T_672 = _T_659[0:0]; // @[LZD.scala 49:47]
  assign _T_673 = _T_666[0:0]; // @[LZD.scala 49:59]
  assign _T_674 = _T_667 ? _T_672 : _T_673; // @[LZD.scala 49:35]
  assign _T_676 = {_T_669,_T_671,_T_674}; // @[Cat.scala 29:58]
  assign _T_677 = _T_651[3:0]; // @[LZD.scala 44:32]
  assign _T_678 = _T_677[3:2]; // @[LZD.scala 43:32]
  assign _T_679 = _T_678 != 2'h0; // @[LZD.scala 39:14]
  assign _T_680 = _T_678[1]; // @[LZD.scala 39:21]
  assign _T_681 = _T_678[0]; // @[LZD.scala 39:30]
  assign _T_682 = ~ _T_681; // @[LZD.scala 39:27]
  assign _T_683 = _T_680 | _T_682; // @[LZD.scala 39:25]
  assign _T_684 = {_T_679,_T_683}; // @[Cat.scala 29:58]
  assign _T_685 = _T_677[1:0]; // @[LZD.scala 44:32]
  assign _T_686 = _T_685 != 2'h0; // @[LZD.scala 39:14]
  assign _T_687 = _T_685[1]; // @[LZD.scala 39:21]
  assign _T_688 = _T_685[0]; // @[LZD.scala 39:30]
  assign _T_689 = ~ _T_688; // @[LZD.scala 39:27]
  assign _T_690 = _T_687 | _T_689; // @[LZD.scala 39:25]
  assign _T_691 = {_T_686,_T_690}; // @[Cat.scala 29:58]
  assign _T_692 = _T_684[1]; // @[Shift.scala 12:21]
  assign _T_693 = _T_691[1]; // @[Shift.scala 12:21]
  assign _T_694 = _T_692 | _T_693; // @[LZD.scala 49:16]
  assign _T_695 = ~ _T_693; // @[LZD.scala 49:27]
  assign _T_696 = _T_692 | _T_695; // @[LZD.scala 49:25]
  assign _T_697 = _T_684[0:0]; // @[LZD.scala 49:47]
  assign _T_698 = _T_691[0:0]; // @[LZD.scala 49:59]
  assign _T_699 = _T_692 ? _T_697 : _T_698; // @[LZD.scala 49:35]
  assign _T_701 = {_T_694,_T_696,_T_699}; // @[Cat.scala 29:58]
  assign _T_702 = _T_676[2]; // @[Shift.scala 12:21]
  assign _T_703 = _T_701[2]; // @[Shift.scala 12:21]
  assign _T_704 = _T_702 | _T_703; // @[LZD.scala 49:16]
  assign _T_705 = ~ _T_703; // @[LZD.scala 49:27]
  assign _T_706 = _T_702 | _T_705; // @[LZD.scala 49:25]
  assign _T_707 = _T_676[1:0]; // @[LZD.scala 49:47]
  assign _T_708 = _T_701[1:0]; // @[LZD.scala 49:59]
  assign _T_709 = _T_702 ? _T_707 : _T_708; // @[LZD.scala 49:35]
  assign _T_711 = {_T_704,_T_706,_T_709}; // @[Cat.scala 29:58]
  assign _T_712 = _T_650[3]; // @[Shift.scala 12:21]
  assign _T_713 = _T_711[3]; // @[Shift.scala 12:21]
  assign _T_714 = _T_712 | _T_713; // @[LZD.scala 49:16]
  assign _T_715 = ~ _T_713; // @[LZD.scala 49:27]
  assign _T_716 = _T_712 | _T_715; // @[LZD.scala 49:25]
  assign _T_717 = _T_650[2:0]; // @[LZD.scala 49:47]
  assign _T_718 = _T_711[2:0]; // @[LZD.scala 49:59]
  assign _T_719 = _T_712 ? _T_717 : _T_718; // @[LZD.scala 49:35]
  assign _T_721 = {_T_714,_T_716,_T_719}; // @[Cat.scala 29:58]
  assign _T_722 = _T_588[10:0]; // @[LZD.scala 44:32]
  assign _T_723 = _T_722[10:3]; // @[LZD.scala 43:32]
  assign _T_724 = _T_723[7:4]; // @[LZD.scala 43:32]
  assign _T_725 = _T_724[3:2]; // @[LZD.scala 43:32]
  assign _T_726 = _T_725 != 2'h0; // @[LZD.scala 39:14]
  assign _T_727 = _T_725[1]; // @[LZD.scala 39:21]
  assign _T_728 = _T_725[0]; // @[LZD.scala 39:30]
  assign _T_729 = ~ _T_728; // @[LZD.scala 39:27]
  assign _T_730 = _T_727 | _T_729; // @[LZD.scala 39:25]
  assign _T_731 = {_T_726,_T_730}; // @[Cat.scala 29:58]
  assign _T_732 = _T_724[1:0]; // @[LZD.scala 44:32]
  assign _T_733 = _T_732 != 2'h0; // @[LZD.scala 39:14]
  assign _T_734 = _T_732[1]; // @[LZD.scala 39:21]
  assign _T_735 = _T_732[0]; // @[LZD.scala 39:30]
  assign _T_736 = ~ _T_735; // @[LZD.scala 39:27]
  assign _T_737 = _T_734 | _T_736; // @[LZD.scala 39:25]
  assign _T_738 = {_T_733,_T_737}; // @[Cat.scala 29:58]
  assign _T_739 = _T_731[1]; // @[Shift.scala 12:21]
  assign _T_740 = _T_738[1]; // @[Shift.scala 12:21]
  assign _T_741 = _T_739 | _T_740; // @[LZD.scala 49:16]
  assign _T_742 = ~ _T_740; // @[LZD.scala 49:27]
  assign _T_743 = _T_739 | _T_742; // @[LZD.scala 49:25]
  assign _T_744 = _T_731[0:0]; // @[LZD.scala 49:47]
  assign _T_745 = _T_738[0:0]; // @[LZD.scala 49:59]
  assign _T_746 = _T_739 ? _T_744 : _T_745; // @[LZD.scala 49:35]
  assign _T_748 = {_T_741,_T_743,_T_746}; // @[Cat.scala 29:58]
  assign _T_749 = _T_723[3:0]; // @[LZD.scala 44:32]
  assign _T_750 = _T_749[3:2]; // @[LZD.scala 43:32]
  assign _T_751 = _T_750 != 2'h0; // @[LZD.scala 39:14]
  assign _T_752 = _T_750[1]; // @[LZD.scala 39:21]
  assign _T_753 = _T_750[0]; // @[LZD.scala 39:30]
  assign _T_754 = ~ _T_753; // @[LZD.scala 39:27]
  assign _T_755 = _T_752 | _T_754; // @[LZD.scala 39:25]
  assign _T_756 = {_T_751,_T_755}; // @[Cat.scala 29:58]
  assign _T_757 = _T_749[1:0]; // @[LZD.scala 44:32]
  assign _T_758 = _T_757 != 2'h0; // @[LZD.scala 39:14]
  assign _T_759 = _T_757[1]; // @[LZD.scala 39:21]
  assign _T_760 = _T_757[0]; // @[LZD.scala 39:30]
  assign _T_761 = ~ _T_760; // @[LZD.scala 39:27]
  assign _T_762 = _T_759 | _T_761; // @[LZD.scala 39:25]
  assign _T_763 = {_T_758,_T_762}; // @[Cat.scala 29:58]
  assign _T_764 = _T_756[1]; // @[Shift.scala 12:21]
  assign _T_765 = _T_763[1]; // @[Shift.scala 12:21]
  assign _T_766 = _T_764 | _T_765; // @[LZD.scala 49:16]
  assign _T_767 = ~ _T_765; // @[LZD.scala 49:27]
  assign _T_768 = _T_764 | _T_767; // @[LZD.scala 49:25]
  assign _T_769 = _T_756[0:0]; // @[LZD.scala 49:47]
  assign _T_770 = _T_763[0:0]; // @[LZD.scala 49:59]
  assign _T_771 = _T_764 ? _T_769 : _T_770; // @[LZD.scala 49:35]
  assign _T_773 = {_T_766,_T_768,_T_771}; // @[Cat.scala 29:58]
  assign _T_774 = _T_748[2]; // @[Shift.scala 12:21]
  assign _T_775 = _T_773[2]; // @[Shift.scala 12:21]
  assign _T_776 = _T_774 | _T_775; // @[LZD.scala 49:16]
  assign _T_777 = ~ _T_775; // @[LZD.scala 49:27]
  assign _T_778 = _T_774 | _T_777; // @[LZD.scala 49:25]
  assign _T_779 = _T_748[1:0]; // @[LZD.scala 49:47]
  assign _T_780 = _T_773[1:0]; // @[LZD.scala 49:59]
  assign _T_781 = _T_774 ? _T_779 : _T_780; // @[LZD.scala 49:35]
  assign _T_783 = {_T_776,_T_778,_T_781}; // @[Cat.scala 29:58]
  assign _T_784 = _T_722[2:0]; // @[LZD.scala 44:32]
  assign _T_785 = _T_784[2:1]; // @[LZD.scala 43:32]
  assign _T_786 = _T_785 != 2'h0; // @[LZD.scala 39:14]
  assign _T_787 = _T_785[1]; // @[LZD.scala 39:21]
  assign _T_788 = _T_785[0]; // @[LZD.scala 39:30]
  assign _T_789 = ~ _T_788; // @[LZD.scala 39:27]
  assign _T_790 = _T_787 | _T_789; // @[LZD.scala 39:25]
  assign _T_791 = {_T_786,_T_790}; // @[Cat.scala 29:58]
  assign _T_792 = _T_784[0:0]; // @[LZD.scala 44:32]
  assign _T_794 = _T_791[1]; // @[Shift.scala 12:21]
  assign _T_796 = _T_791[0:0]; // @[LZD.scala 55:32]
  assign _T_797 = _T_794 ? _T_796 : _T_792; // @[LZD.scala 55:20]
  assign _T_799 = _T_783[3]; // @[Shift.scala 12:21]
  assign _T_801 = {1'h1,_T_794,_T_797}; // @[Cat.scala 29:58]
  assign _T_802 = _T_783[2:0]; // @[LZD.scala 55:32]
  assign _T_803 = _T_799 ? _T_802 : _T_801; // @[LZD.scala 55:20]
  assign _T_804 = {_T_799,_T_803}; // @[Cat.scala 29:58]
  assign _T_805 = _T_721[4]; // @[Shift.scala 12:21]
  assign _T_807 = _T_721[3:0]; // @[LZD.scala 55:32]
  assign _T_808 = _T_805 ? _T_807 : _T_804; // @[LZD.scala 55:20]
  assign _T_809 = {_T_805,_T_808}; // @[Cat.scala 29:58]
  assign _T_810 = ~ _T_809; // @[convert.scala 21:22]
  assign _T_811 = realC[25:0]; // @[convert.scala 22:36]
  assign _T_812 = _T_810 < 5'h1a; // @[Shift.scala 16:24]
  assign _T_814 = _T_810[4]; // @[Shift.scala 12:21]
  assign _T_815 = _T_811[9:0]; // @[Shift.scala 64:52]
  assign _T_817 = {_T_815,16'h0}; // @[Cat.scala 29:58]
  assign _T_818 = _T_814 ? _T_817 : _T_811; // @[Shift.scala 64:27]
  assign _T_819 = _T_810[3:0]; // @[Shift.scala 66:70]
  assign _T_820 = _T_819[3]; // @[Shift.scala 12:21]
  assign _T_821 = _T_818[17:0]; // @[Shift.scala 64:52]
  assign _T_823 = {_T_821,8'h0}; // @[Cat.scala 29:58]
  assign _T_824 = _T_820 ? _T_823 : _T_818; // @[Shift.scala 64:27]
  assign _T_825 = _T_819[2:0]; // @[Shift.scala 66:70]
  assign _T_826 = _T_825[2]; // @[Shift.scala 12:21]
  assign _T_827 = _T_824[21:0]; // @[Shift.scala 64:52]
  assign _T_829 = {_T_827,4'h0}; // @[Cat.scala 29:58]
  assign _T_830 = _T_826 ? _T_829 : _T_824; // @[Shift.scala 64:27]
  assign _T_831 = _T_825[1:0]; // @[Shift.scala 66:70]
  assign _T_832 = _T_831[1]; // @[Shift.scala 12:21]
  assign _T_833 = _T_830[23:0]; // @[Shift.scala 64:52]
  assign _T_835 = {_T_833,2'h0}; // @[Cat.scala 29:58]
  assign _T_836 = _T_832 ? _T_835 : _T_830; // @[Shift.scala 64:27]
  assign _T_837 = _T_831[0:0]; // @[Shift.scala 66:70]
  assign _T_839 = _T_836[24:0]; // @[Shift.scala 64:52]
  assign _T_840 = {_T_839,1'h0}; // @[Cat.scala 29:58]
  assign _T_841 = _T_837 ? _T_840 : _T_836; // @[Shift.scala 64:27]
  assign _T_842 = _T_812 ? _T_841 : 26'h0; // @[Shift.scala 16:10]
  assign _T_843 = _T_842[25:23]; // @[convert.scala 23:34]
  assign decC_fraction = _T_842[22:0]; // @[convert.scala 24:34]
  assign _T_845 = _T_585 == 1'h0; // @[convert.scala 25:26]
  assign _T_847 = _T_585 ? _T_810 : _T_809; // @[convert.scala 25:42]
  assign _T_850 = ~ _T_843; // @[convert.scala 26:67]
  assign _T_851 = _T_583 ? _T_850 : _T_843; // @[convert.scala 26:51]
  assign _T_852 = {_T_845,_T_847,_T_851}; // @[Cat.scala 29:58]
  assign _T_854 = realC[27:0]; // @[convert.scala 29:56]
  assign _T_855 = _T_854 != 28'h0; // @[convert.scala 29:60]
  assign _T_856 = ~ _T_855; // @[convert.scala 29:41]
  assign decC_isNaR = _T_583 & _T_856; // @[convert.scala 29:39]
  assign _T_859 = _T_583 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_859 & _T_856; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_852); // @[convert.scala 32:24]
  assign _T_867 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_867 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_868 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_869 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_870 = _T_868 & _T_869; // @[PositFMA.scala 59:45]
  assign _T_872 = {_T_13,_T_870,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_872); // @[PositFMA.scala 59:76]
  assign _T_873 = ~ _T_298; // @[PositFMA.scala 60:34]
  assign _T_874 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_875 = _T_873 & _T_874; // @[PositFMA.scala 60:45]
  assign _T_877 = {_T_298,_T_875,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_877); // @[PositFMA.scala 60:76]
  assign _T_878 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_878); // @[PositFMA.scala 61:33]
  assign _T_879 = sigP[46:0]; // @[PositFMA.scala 62:29]
  assign _T_880 = _T_879 != 47'h0; // @[PositFMA.scala 62:33]
  assign eqTwo = ~ _T_880; // @[PositFMA.scala 62:19]
  assign _T_881 = sigP[48]; // @[PositFMA.scala 64:29]
  assign _T_882 = sigP[47]; // @[PositFMA.scala 64:56]
  assign _T_883 = ~ _T_882; // @[PositFMA.scala 64:51]
  assign _T_884 = _T_881 & _T_883; // @[PositFMA.scala 64:49]
  assign eqFour = _T_884 & eqTwo; // @[PositFMA.scala 64:76]
  assign _T_885 = sigP[49]; // @[PositFMA.scala 66:23]
  assign geTwo = _T_885 ^ _T_882; // @[PositFMA.scala 66:43]
  assign _T_887 = {eqFour,geTwo}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_887)}; // @[PositFMA.scala 67:38]
  assign mulSign = sigP[49:49]; // @[PositFMA.scala 68:28]
  assign _T_888 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 70:30]
  assign _GEN_12 = {{7{expBias[2]}},expBias}; // @[PositFMA.scala 70:44]
  assign _T_890 = $signed(_T_888) + $signed(_GEN_12); // @[PositFMA.scala 70:44]
  assign mulScale = $signed(_T_890); // @[PositFMA.scala 70:44]
  assign _T_891 = sigP[47:0]; // @[PositFMA.scala 73:29]
  assign _T_892 = sigP[46:0]; // @[PositFMA.scala 74:29]
  assign _T_893 = {_T_892, 1'h0}; // @[PositFMA.scala 74:48]
  assign mulSigTmp = geTwo ? _T_891 : _T_893; // @[PositFMA.scala 71:22]
  assign _T_895 = mulSigTmp[47:47]; // @[PositFMA.scala 78:39]
  assign _T_896 = _T_895 | eqFour; // @[PositFMA.scala 78:43]
  assign _T_897 = mulSigTmp[46:0]; // @[PositFMA.scala 79:39]
  assign mulSig = {mulSign,_T_896,_T_897}; // @[Cat.scala 29:58]
  assign _T_923 = ~ addSign_phase2; // @[PositFMA.scala 108:29]
  assign _T_924 = ~ addZero_phase2; // @[PositFMA.scala 108:47]
  assign _T_925 = _T_923 & _T_924; // @[PositFMA.scala 108:45]
  assign extAddSig = {addSign_phase2,_T_925,addFrac_phase2,24'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[8]}},addScale_phase2}; // @[PositFMA.scala 112:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 112:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[8]}},addScale_phase2}); // @[PositFMA.scala 113:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[8]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 114:26]
  assign _T_929 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 115:36]
  assign scaleDiff = $signed(_T_929); // @[PositFMA.scala 115:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 116:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 117:26]
  assign _T_930 = $unsigned(scaleDiff); // @[PositFMA.scala 118:69]
  assign _T_931 = _T_930 < 10'h31; // @[Shift.scala 39:24]
  assign _T_932 = _T_930[5:0]; // @[Shift.scala 40:44]
  assign _T_933 = smallerSigTmp[48:32]; // @[Shift.scala 90:30]
  assign _T_934 = smallerSigTmp[31:0]; // @[Shift.scala 90:48]
  assign _T_935 = _T_934 != 32'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{16'd0}, _T_935}; // @[Shift.scala 90:39]
  assign _T_936 = _T_933 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_937 = _T_932[5]; // @[Shift.scala 12:21]
  assign _T_938 = smallerSigTmp[48]; // @[Shift.scala 12:21]
  assign _T_940 = _T_938 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_941 = {_T_940,_T_936}; // @[Cat.scala 29:58]
  assign _T_942 = _T_937 ? _T_941 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_943 = _T_932[4:0]; // @[Shift.scala 92:77]
  assign _T_944 = _T_942[48:16]; // @[Shift.scala 90:30]
  assign _T_945 = _T_942[15:0]; // @[Shift.scala 90:48]
  assign _T_946 = _T_945 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{32'd0}, _T_946}; // @[Shift.scala 90:39]
  assign _T_947 = _T_944 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_948 = _T_943[4]; // @[Shift.scala 12:21]
  assign _T_949 = _T_942[48]; // @[Shift.scala 12:21]
  assign _T_951 = _T_949 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_952 = {_T_951,_T_947}; // @[Cat.scala 29:58]
  assign _T_953 = _T_948 ? _T_952 : _T_942; // @[Shift.scala 91:22]
  assign _T_954 = _T_943[3:0]; // @[Shift.scala 92:77]
  assign _T_955 = _T_953[48:8]; // @[Shift.scala 90:30]
  assign _T_956 = _T_953[7:0]; // @[Shift.scala 90:48]
  assign _T_957 = _T_956 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{40'd0}, _T_957}; // @[Shift.scala 90:39]
  assign _T_958 = _T_955 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_959 = _T_954[3]; // @[Shift.scala 12:21]
  assign _T_960 = _T_953[48]; // @[Shift.scala 12:21]
  assign _T_962 = _T_960 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_963 = {_T_962,_T_958}; // @[Cat.scala 29:58]
  assign _T_964 = _T_959 ? _T_963 : _T_953; // @[Shift.scala 91:22]
  assign _T_965 = _T_954[2:0]; // @[Shift.scala 92:77]
  assign _T_966 = _T_964[48:4]; // @[Shift.scala 90:30]
  assign _T_967 = _T_964[3:0]; // @[Shift.scala 90:48]
  assign _T_968 = _T_967 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_17 = {{44'd0}, _T_968}; // @[Shift.scala 90:39]
  assign _T_969 = _T_966 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_970 = _T_965[2]; // @[Shift.scala 12:21]
  assign _T_971 = _T_964[48]; // @[Shift.scala 12:21]
  assign _T_973 = _T_971 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_974 = {_T_973,_T_969}; // @[Cat.scala 29:58]
  assign _T_975 = _T_970 ? _T_974 : _T_964; // @[Shift.scala 91:22]
  assign _T_976 = _T_965[1:0]; // @[Shift.scala 92:77]
  assign _T_977 = _T_975[48:2]; // @[Shift.scala 90:30]
  assign _T_978 = _T_975[1:0]; // @[Shift.scala 90:48]
  assign _T_979 = _T_978 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_18 = {{46'd0}, _T_979}; // @[Shift.scala 90:39]
  assign _T_980 = _T_977 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_981 = _T_976[1]; // @[Shift.scala 12:21]
  assign _T_982 = _T_975[48]; // @[Shift.scala 12:21]
  assign _T_984 = _T_982 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_985 = {_T_984,_T_980}; // @[Cat.scala 29:58]
  assign _T_986 = _T_981 ? _T_985 : _T_975; // @[Shift.scala 91:22]
  assign _T_987 = _T_976[0:0]; // @[Shift.scala 92:77]
  assign _T_988 = _T_986[48:1]; // @[Shift.scala 90:30]
  assign _T_989 = _T_986[0:0]; // @[Shift.scala 90:48]
  assign _GEN_19 = {{47'd0}, _T_989}; // @[Shift.scala 90:39]
  assign _T_991 = _T_988 | _GEN_19; // @[Shift.scala 90:39]
  assign _T_993 = _T_986[48]; // @[Shift.scala 12:21]
  assign _T_994 = {_T_993,_T_991}; // @[Cat.scala 29:58]
  assign _T_995 = _T_987 ? _T_994 : _T_986; // @[Shift.scala 91:22]
  assign _T_998 = _T_938 ? 49'h1ffffffffffff : 49'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_931 ? _T_995 : _T_998; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 119:34]
  assign _T_999 = mulSig_phase2[48:48]; // @[PositFMA.scala 120:42]
  assign _T_1000 = _T_999 ^ addSign_phase2; // @[PositFMA.scala 120:46]
  assign _T_1001 = rawSumSig[49:49]; // @[PositFMA.scala 120:79]
  assign sumSign = _T_1000 ^ _T_1001; // @[PositFMA.scala 120:63]
  assign _T_1003 = greaterSig + smallerSig; // @[PositFMA.scala 121:50]
  assign signSumSig = {sumSign,_T_1003}; // @[Cat.scala 29:58]
  assign _T_1004 = signSumSig[49:1]; // @[PositFMA.scala 125:33]
  assign _T_1005 = signSumSig[48:0]; // @[PositFMA.scala 125:68]
  assign sumXor = _T_1004 ^ _T_1005; // @[PositFMA.scala 125:51]
  assign _T_1006 = sumXor[48:17]; // @[LZD.scala 43:32]
  assign _T_1007 = _T_1006[31:16]; // @[LZD.scala 43:32]
  assign _T_1008 = _T_1007[15:8]; // @[LZD.scala 43:32]
  assign _T_1009 = _T_1008[7:4]; // @[LZD.scala 43:32]
  assign _T_1010 = _T_1009[3:2]; // @[LZD.scala 43:32]
  assign _T_1011 = _T_1010 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1012 = _T_1010[1]; // @[LZD.scala 39:21]
  assign _T_1013 = _T_1010[0]; // @[LZD.scala 39:30]
  assign _T_1014 = ~ _T_1013; // @[LZD.scala 39:27]
  assign _T_1015 = _T_1012 | _T_1014; // @[LZD.scala 39:25]
  assign _T_1016 = {_T_1011,_T_1015}; // @[Cat.scala 29:58]
  assign _T_1017 = _T_1009[1:0]; // @[LZD.scala 44:32]
  assign _T_1018 = _T_1017 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1019 = _T_1017[1]; // @[LZD.scala 39:21]
  assign _T_1020 = _T_1017[0]; // @[LZD.scala 39:30]
  assign _T_1021 = ~ _T_1020; // @[LZD.scala 39:27]
  assign _T_1022 = _T_1019 | _T_1021; // @[LZD.scala 39:25]
  assign _T_1023 = {_T_1018,_T_1022}; // @[Cat.scala 29:58]
  assign _T_1024 = _T_1016[1]; // @[Shift.scala 12:21]
  assign _T_1025 = _T_1023[1]; // @[Shift.scala 12:21]
  assign _T_1026 = _T_1024 | _T_1025; // @[LZD.scala 49:16]
  assign _T_1027 = ~ _T_1025; // @[LZD.scala 49:27]
  assign _T_1028 = _T_1024 | _T_1027; // @[LZD.scala 49:25]
  assign _T_1029 = _T_1016[0:0]; // @[LZD.scala 49:47]
  assign _T_1030 = _T_1023[0:0]; // @[LZD.scala 49:59]
  assign _T_1031 = _T_1024 ? _T_1029 : _T_1030; // @[LZD.scala 49:35]
  assign _T_1033 = {_T_1026,_T_1028,_T_1031}; // @[Cat.scala 29:58]
  assign _T_1034 = _T_1008[3:0]; // @[LZD.scala 44:32]
  assign _T_1035 = _T_1034[3:2]; // @[LZD.scala 43:32]
  assign _T_1036 = _T_1035 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1037 = _T_1035[1]; // @[LZD.scala 39:21]
  assign _T_1038 = _T_1035[0]; // @[LZD.scala 39:30]
  assign _T_1039 = ~ _T_1038; // @[LZD.scala 39:27]
  assign _T_1040 = _T_1037 | _T_1039; // @[LZD.scala 39:25]
  assign _T_1041 = {_T_1036,_T_1040}; // @[Cat.scala 29:58]
  assign _T_1042 = _T_1034[1:0]; // @[LZD.scala 44:32]
  assign _T_1043 = _T_1042 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1044 = _T_1042[1]; // @[LZD.scala 39:21]
  assign _T_1045 = _T_1042[0]; // @[LZD.scala 39:30]
  assign _T_1046 = ~ _T_1045; // @[LZD.scala 39:27]
  assign _T_1047 = _T_1044 | _T_1046; // @[LZD.scala 39:25]
  assign _T_1048 = {_T_1043,_T_1047}; // @[Cat.scala 29:58]
  assign _T_1049 = _T_1041[1]; // @[Shift.scala 12:21]
  assign _T_1050 = _T_1048[1]; // @[Shift.scala 12:21]
  assign _T_1051 = _T_1049 | _T_1050; // @[LZD.scala 49:16]
  assign _T_1052 = ~ _T_1050; // @[LZD.scala 49:27]
  assign _T_1053 = _T_1049 | _T_1052; // @[LZD.scala 49:25]
  assign _T_1054 = _T_1041[0:0]; // @[LZD.scala 49:47]
  assign _T_1055 = _T_1048[0:0]; // @[LZD.scala 49:59]
  assign _T_1056 = _T_1049 ? _T_1054 : _T_1055; // @[LZD.scala 49:35]
  assign _T_1058 = {_T_1051,_T_1053,_T_1056}; // @[Cat.scala 29:58]
  assign _T_1059 = _T_1033[2]; // @[Shift.scala 12:21]
  assign _T_1060 = _T_1058[2]; // @[Shift.scala 12:21]
  assign _T_1061 = _T_1059 | _T_1060; // @[LZD.scala 49:16]
  assign _T_1062 = ~ _T_1060; // @[LZD.scala 49:27]
  assign _T_1063 = _T_1059 | _T_1062; // @[LZD.scala 49:25]
  assign _T_1064 = _T_1033[1:0]; // @[LZD.scala 49:47]
  assign _T_1065 = _T_1058[1:0]; // @[LZD.scala 49:59]
  assign _T_1066 = _T_1059 ? _T_1064 : _T_1065; // @[LZD.scala 49:35]
  assign _T_1068 = {_T_1061,_T_1063,_T_1066}; // @[Cat.scala 29:58]
  assign _T_1069 = _T_1007[7:0]; // @[LZD.scala 44:32]
  assign _T_1070 = _T_1069[7:4]; // @[LZD.scala 43:32]
  assign _T_1071 = _T_1070[3:2]; // @[LZD.scala 43:32]
  assign _T_1072 = _T_1071 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1073 = _T_1071[1]; // @[LZD.scala 39:21]
  assign _T_1074 = _T_1071[0]; // @[LZD.scala 39:30]
  assign _T_1075 = ~ _T_1074; // @[LZD.scala 39:27]
  assign _T_1076 = _T_1073 | _T_1075; // @[LZD.scala 39:25]
  assign _T_1077 = {_T_1072,_T_1076}; // @[Cat.scala 29:58]
  assign _T_1078 = _T_1070[1:0]; // @[LZD.scala 44:32]
  assign _T_1079 = _T_1078 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1080 = _T_1078[1]; // @[LZD.scala 39:21]
  assign _T_1081 = _T_1078[0]; // @[LZD.scala 39:30]
  assign _T_1082 = ~ _T_1081; // @[LZD.scala 39:27]
  assign _T_1083 = _T_1080 | _T_1082; // @[LZD.scala 39:25]
  assign _T_1084 = {_T_1079,_T_1083}; // @[Cat.scala 29:58]
  assign _T_1085 = _T_1077[1]; // @[Shift.scala 12:21]
  assign _T_1086 = _T_1084[1]; // @[Shift.scala 12:21]
  assign _T_1087 = _T_1085 | _T_1086; // @[LZD.scala 49:16]
  assign _T_1088 = ~ _T_1086; // @[LZD.scala 49:27]
  assign _T_1089 = _T_1085 | _T_1088; // @[LZD.scala 49:25]
  assign _T_1090 = _T_1077[0:0]; // @[LZD.scala 49:47]
  assign _T_1091 = _T_1084[0:0]; // @[LZD.scala 49:59]
  assign _T_1092 = _T_1085 ? _T_1090 : _T_1091; // @[LZD.scala 49:35]
  assign _T_1094 = {_T_1087,_T_1089,_T_1092}; // @[Cat.scala 29:58]
  assign _T_1095 = _T_1069[3:0]; // @[LZD.scala 44:32]
  assign _T_1096 = _T_1095[3:2]; // @[LZD.scala 43:32]
  assign _T_1097 = _T_1096 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1098 = _T_1096[1]; // @[LZD.scala 39:21]
  assign _T_1099 = _T_1096[0]; // @[LZD.scala 39:30]
  assign _T_1100 = ~ _T_1099; // @[LZD.scala 39:27]
  assign _T_1101 = _T_1098 | _T_1100; // @[LZD.scala 39:25]
  assign _T_1102 = {_T_1097,_T_1101}; // @[Cat.scala 29:58]
  assign _T_1103 = _T_1095[1:0]; // @[LZD.scala 44:32]
  assign _T_1104 = _T_1103 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1105 = _T_1103[1]; // @[LZD.scala 39:21]
  assign _T_1106 = _T_1103[0]; // @[LZD.scala 39:30]
  assign _T_1107 = ~ _T_1106; // @[LZD.scala 39:27]
  assign _T_1108 = _T_1105 | _T_1107; // @[LZD.scala 39:25]
  assign _T_1109 = {_T_1104,_T_1108}; // @[Cat.scala 29:58]
  assign _T_1110 = _T_1102[1]; // @[Shift.scala 12:21]
  assign _T_1111 = _T_1109[1]; // @[Shift.scala 12:21]
  assign _T_1112 = _T_1110 | _T_1111; // @[LZD.scala 49:16]
  assign _T_1113 = ~ _T_1111; // @[LZD.scala 49:27]
  assign _T_1114 = _T_1110 | _T_1113; // @[LZD.scala 49:25]
  assign _T_1115 = _T_1102[0:0]; // @[LZD.scala 49:47]
  assign _T_1116 = _T_1109[0:0]; // @[LZD.scala 49:59]
  assign _T_1117 = _T_1110 ? _T_1115 : _T_1116; // @[LZD.scala 49:35]
  assign _T_1119 = {_T_1112,_T_1114,_T_1117}; // @[Cat.scala 29:58]
  assign _T_1120 = _T_1094[2]; // @[Shift.scala 12:21]
  assign _T_1121 = _T_1119[2]; // @[Shift.scala 12:21]
  assign _T_1122 = _T_1120 | _T_1121; // @[LZD.scala 49:16]
  assign _T_1123 = ~ _T_1121; // @[LZD.scala 49:27]
  assign _T_1124 = _T_1120 | _T_1123; // @[LZD.scala 49:25]
  assign _T_1125 = _T_1094[1:0]; // @[LZD.scala 49:47]
  assign _T_1126 = _T_1119[1:0]; // @[LZD.scala 49:59]
  assign _T_1127 = _T_1120 ? _T_1125 : _T_1126; // @[LZD.scala 49:35]
  assign _T_1129 = {_T_1122,_T_1124,_T_1127}; // @[Cat.scala 29:58]
  assign _T_1130 = _T_1068[3]; // @[Shift.scala 12:21]
  assign _T_1131 = _T_1129[3]; // @[Shift.scala 12:21]
  assign _T_1132 = _T_1130 | _T_1131; // @[LZD.scala 49:16]
  assign _T_1133 = ~ _T_1131; // @[LZD.scala 49:27]
  assign _T_1134 = _T_1130 | _T_1133; // @[LZD.scala 49:25]
  assign _T_1135 = _T_1068[2:0]; // @[LZD.scala 49:47]
  assign _T_1136 = _T_1129[2:0]; // @[LZD.scala 49:59]
  assign _T_1137 = _T_1130 ? _T_1135 : _T_1136; // @[LZD.scala 49:35]
  assign _T_1139 = {_T_1132,_T_1134,_T_1137}; // @[Cat.scala 29:58]
  assign _T_1140 = _T_1006[15:0]; // @[LZD.scala 44:32]
  assign _T_1141 = _T_1140[15:8]; // @[LZD.scala 43:32]
  assign _T_1142 = _T_1141[7:4]; // @[LZD.scala 43:32]
  assign _T_1143 = _T_1142[3:2]; // @[LZD.scala 43:32]
  assign _T_1144 = _T_1143 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1145 = _T_1143[1]; // @[LZD.scala 39:21]
  assign _T_1146 = _T_1143[0]; // @[LZD.scala 39:30]
  assign _T_1147 = ~ _T_1146; // @[LZD.scala 39:27]
  assign _T_1148 = _T_1145 | _T_1147; // @[LZD.scala 39:25]
  assign _T_1149 = {_T_1144,_T_1148}; // @[Cat.scala 29:58]
  assign _T_1150 = _T_1142[1:0]; // @[LZD.scala 44:32]
  assign _T_1151 = _T_1150 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1152 = _T_1150[1]; // @[LZD.scala 39:21]
  assign _T_1153 = _T_1150[0]; // @[LZD.scala 39:30]
  assign _T_1154 = ~ _T_1153; // @[LZD.scala 39:27]
  assign _T_1155 = _T_1152 | _T_1154; // @[LZD.scala 39:25]
  assign _T_1156 = {_T_1151,_T_1155}; // @[Cat.scala 29:58]
  assign _T_1157 = _T_1149[1]; // @[Shift.scala 12:21]
  assign _T_1158 = _T_1156[1]; // @[Shift.scala 12:21]
  assign _T_1159 = _T_1157 | _T_1158; // @[LZD.scala 49:16]
  assign _T_1160 = ~ _T_1158; // @[LZD.scala 49:27]
  assign _T_1161 = _T_1157 | _T_1160; // @[LZD.scala 49:25]
  assign _T_1162 = _T_1149[0:0]; // @[LZD.scala 49:47]
  assign _T_1163 = _T_1156[0:0]; // @[LZD.scala 49:59]
  assign _T_1164 = _T_1157 ? _T_1162 : _T_1163; // @[LZD.scala 49:35]
  assign _T_1166 = {_T_1159,_T_1161,_T_1164}; // @[Cat.scala 29:58]
  assign _T_1167 = _T_1141[3:0]; // @[LZD.scala 44:32]
  assign _T_1168 = _T_1167[3:2]; // @[LZD.scala 43:32]
  assign _T_1169 = _T_1168 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1170 = _T_1168[1]; // @[LZD.scala 39:21]
  assign _T_1171 = _T_1168[0]; // @[LZD.scala 39:30]
  assign _T_1172 = ~ _T_1171; // @[LZD.scala 39:27]
  assign _T_1173 = _T_1170 | _T_1172; // @[LZD.scala 39:25]
  assign _T_1174 = {_T_1169,_T_1173}; // @[Cat.scala 29:58]
  assign _T_1175 = _T_1167[1:0]; // @[LZD.scala 44:32]
  assign _T_1176 = _T_1175 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1177 = _T_1175[1]; // @[LZD.scala 39:21]
  assign _T_1178 = _T_1175[0]; // @[LZD.scala 39:30]
  assign _T_1179 = ~ _T_1178; // @[LZD.scala 39:27]
  assign _T_1180 = _T_1177 | _T_1179; // @[LZD.scala 39:25]
  assign _T_1181 = {_T_1176,_T_1180}; // @[Cat.scala 29:58]
  assign _T_1182 = _T_1174[1]; // @[Shift.scala 12:21]
  assign _T_1183 = _T_1181[1]; // @[Shift.scala 12:21]
  assign _T_1184 = _T_1182 | _T_1183; // @[LZD.scala 49:16]
  assign _T_1185 = ~ _T_1183; // @[LZD.scala 49:27]
  assign _T_1186 = _T_1182 | _T_1185; // @[LZD.scala 49:25]
  assign _T_1187 = _T_1174[0:0]; // @[LZD.scala 49:47]
  assign _T_1188 = _T_1181[0:0]; // @[LZD.scala 49:59]
  assign _T_1189 = _T_1182 ? _T_1187 : _T_1188; // @[LZD.scala 49:35]
  assign _T_1191 = {_T_1184,_T_1186,_T_1189}; // @[Cat.scala 29:58]
  assign _T_1192 = _T_1166[2]; // @[Shift.scala 12:21]
  assign _T_1193 = _T_1191[2]; // @[Shift.scala 12:21]
  assign _T_1194 = _T_1192 | _T_1193; // @[LZD.scala 49:16]
  assign _T_1195 = ~ _T_1193; // @[LZD.scala 49:27]
  assign _T_1196 = _T_1192 | _T_1195; // @[LZD.scala 49:25]
  assign _T_1197 = _T_1166[1:0]; // @[LZD.scala 49:47]
  assign _T_1198 = _T_1191[1:0]; // @[LZD.scala 49:59]
  assign _T_1199 = _T_1192 ? _T_1197 : _T_1198; // @[LZD.scala 49:35]
  assign _T_1201 = {_T_1194,_T_1196,_T_1199}; // @[Cat.scala 29:58]
  assign _T_1202 = _T_1140[7:0]; // @[LZD.scala 44:32]
  assign _T_1203 = _T_1202[7:4]; // @[LZD.scala 43:32]
  assign _T_1204 = _T_1203[3:2]; // @[LZD.scala 43:32]
  assign _T_1205 = _T_1204 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1206 = _T_1204[1]; // @[LZD.scala 39:21]
  assign _T_1207 = _T_1204[0]; // @[LZD.scala 39:30]
  assign _T_1208 = ~ _T_1207; // @[LZD.scala 39:27]
  assign _T_1209 = _T_1206 | _T_1208; // @[LZD.scala 39:25]
  assign _T_1210 = {_T_1205,_T_1209}; // @[Cat.scala 29:58]
  assign _T_1211 = _T_1203[1:0]; // @[LZD.scala 44:32]
  assign _T_1212 = _T_1211 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1213 = _T_1211[1]; // @[LZD.scala 39:21]
  assign _T_1214 = _T_1211[0]; // @[LZD.scala 39:30]
  assign _T_1215 = ~ _T_1214; // @[LZD.scala 39:27]
  assign _T_1216 = _T_1213 | _T_1215; // @[LZD.scala 39:25]
  assign _T_1217 = {_T_1212,_T_1216}; // @[Cat.scala 29:58]
  assign _T_1218 = _T_1210[1]; // @[Shift.scala 12:21]
  assign _T_1219 = _T_1217[1]; // @[Shift.scala 12:21]
  assign _T_1220 = _T_1218 | _T_1219; // @[LZD.scala 49:16]
  assign _T_1221 = ~ _T_1219; // @[LZD.scala 49:27]
  assign _T_1222 = _T_1218 | _T_1221; // @[LZD.scala 49:25]
  assign _T_1223 = _T_1210[0:0]; // @[LZD.scala 49:47]
  assign _T_1224 = _T_1217[0:0]; // @[LZD.scala 49:59]
  assign _T_1225 = _T_1218 ? _T_1223 : _T_1224; // @[LZD.scala 49:35]
  assign _T_1227 = {_T_1220,_T_1222,_T_1225}; // @[Cat.scala 29:58]
  assign _T_1228 = _T_1202[3:0]; // @[LZD.scala 44:32]
  assign _T_1229 = _T_1228[3:2]; // @[LZD.scala 43:32]
  assign _T_1230 = _T_1229 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1231 = _T_1229[1]; // @[LZD.scala 39:21]
  assign _T_1232 = _T_1229[0]; // @[LZD.scala 39:30]
  assign _T_1233 = ~ _T_1232; // @[LZD.scala 39:27]
  assign _T_1234 = _T_1231 | _T_1233; // @[LZD.scala 39:25]
  assign _T_1235 = {_T_1230,_T_1234}; // @[Cat.scala 29:58]
  assign _T_1236 = _T_1228[1:0]; // @[LZD.scala 44:32]
  assign _T_1237 = _T_1236 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1238 = _T_1236[1]; // @[LZD.scala 39:21]
  assign _T_1239 = _T_1236[0]; // @[LZD.scala 39:30]
  assign _T_1240 = ~ _T_1239; // @[LZD.scala 39:27]
  assign _T_1241 = _T_1238 | _T_1240; // @[LZD.scala 39:25]
  assign _T_1242 = {_T_1237,_T_1241}; // @[Cat.scala 29:58]
  assign _T_1243 = _T_1235[1]; // @[Shift.scala 12:21]
  assign _T_1244 = _T_1242[1]; // @[Shift.scala 12:21]
  assign _T_1245 = _T_1243 | _T_1244; // @[LZD.scala 49:16]
  assign _T_1246 = ~ _T_1244; // @[LZD.scala 49:27]
  assign _T_1247 = _T_1243 | _T_1246; // @[LZD.scala 49:25]
  assign _T_1248 = _T_1235[0:0]; // @[LZD.scala 49:47]
  assign _T_1249 = _T_1242[0:0]; // @[LZD.scala 49:59]
  assign _T_1250 = _T_1243 ? _T_1248 : _T_1249; // @[LZD.scala 49:35]
  assign _T_1252 = {_T_1245,_T_1247,_T_1250}; // @[Cat.scala 29:58]
  assign _T_1253 = _T_1227[2]; // @[Shift.scala 12:21]
  assign _T_1254 = _T_1252[2]; // @[Shift.scala 12:21]
  assign _T_1255 = _T_1253 | _T_1254; // @[LZD.scala 49:16]
  assign _T_1256 = ~ _T_1254; // @[LZD.scala 49:27]
  assign _T_1257 = _T_1253 | _T_1256; // @[LZD.scala 49:25]
  assign _T_1258 = _T_1227[1:0]; // @[LZD.scala 49:47]
  assign _T_1259 = _T_1252[1:0]; // @[LZD.scala 49:59]
  assign _T_1260 = _T_1253 ? _T_1258 : _T_1259; // @[LZD.scala 49:35]
  assign _T_1262 = {_T_1255,_T_1257,_T_1260}; // @[Cat.scala 29:58]
  assign _T_1263 = _T_1201[3]; // @[Shift.scala 12:21]
  assign _T_1264 = _T_1262[3]; // @[Shift.scala 12:21]
  assign _T_1265 = _T_1263 | _T_1264; // @[LZD.scala 49:16]
  assign _T_1266 = ~ _T_1264; // @[LZD.scala 49:27]
  assign _T_1267 = _T_1263 | _T_1266; // @[LZD.scala 49:25]
  assign _T_1268 = _T_1201[2:0]; // @[LZD.scala 49:47]
  assign _T_1269 = _T_1262[2:0]; // @[LZD.scala 49:59]
  assign _T_1270 = _T_1263 ? _T_1268 : _T_1269; // @[LZD.scala 49:35]
  assign _T_1272 = {_T_1265,_T_1267,_T_1270}; // @[Cat.scala 29:58]
  assign _T_1273 = _T_1139[4]; // @[Shift.scala 12:21]
  assign _T_1274 = _T_1272[4]; // @[Shift.scala 12:21]
  assign _T_1275 = _T_1273 | _T_1274; // @[LZD.scala 49:16]
  assign _T_1276 = ~ _T_1274; // @[LZD.scala 49:27]
  assign _T_1277 = _T_1273 | _T_1276; // @[LZD.scala 49:25]
  assign _T_1278 = _T_1139[3:0]; // @[LZD.scala 49:47]
  assign _T_1279 = _T_1272[3:0]; // @[LZD.scala 49:59]
  assign _T_1280 = _T_1273 ? _T_1278 : _T_1279; // @[LZD.scala 49:35]
  assign _T_1282 = {_T_1275,_T_1277,_T_1280}; // @[Cat.scala 29:58]
  assign _T_1283 = sumXor[16:0]; // @[LZD.scala 44:32]
  assign _T_1284 = _T_1283[16:1]; // @[LZD.scala 43:32]
  assign _T_1285 = _T_1284[15:8]; // @[LZD.scala 43:32]
  assign _T_1286 = _T_1285[7:4]; // @[LZD.scala 43:32]
  assign _T_1287 = _T_1286[3:2]; // @[LZD.scala 43:32]
  assign _T_1288 = _T_1287 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1289 = _T_1287[1]; // @[LZD.scala 39:21]
  assign _T_1290 = _T_1287[0]; // @[LZD.scala 39:30]
  assign _T_1291 = ~ _T_1290; // @[LZD.scala 39:27]
  assign _T_1292 = _T_1289 | _T_1291; // @[LZD.scala 39:25]
  assign _T_1293 = {_T_1288,_T_1292}; // @[Cat.scala 29:58]
  assign _T_1294 = _T_1286[1:0]; // @[LZD.scala 44:32]
  assign _T_1295 = _T_1294 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1296 = _T_1294[1]; // @[LZD.scala 39:21]
  assign _T_1297 = _T_1294[0]; // @[LZD.scala 39:30]
  assign _T_1298 = ~ _T_1297; // @[LZD.scala 39:27]
  assign _T_1299 = _T_1296 | _T_1298; // @[LZD.scala 39:25]
  assign _T_1300 = {_T_1295,_T_1299}; // @[Cat.scala 29:58]
  assign _T_1301 = _T_1293[1]; // @[Shift.scala 12:21]
  assign _T_1302 = _T_1300[1]; // @[Shift.scala 12:21]
  assign _T_1303 = _T_1301 | _T_1302; // @[LZD.scala 49:16]
  assign _T_1304 = ~ _T_1302; // @[LZD.scala 49:27]
  assign _T_1305 = _T_1301 | _T_1304; // @[LZD.scala 49:25]
  assign _T_1306 = _T_1293[0:0]; // @[LZD.scala 49:47]
  assign _T_1307 = _T_1300[0:0]; // @[LZD.scala 49:59]
  assign _T_1308 = _T_1301 ? _T_1306 : _T_1307; // @[LZD.scala 49:35]
  assign _T_1310 = {_T_1303,_T_1305,_T_1308}; // @[Cat.scala 29:58]
  assign _T_1311 = _T_1285[3:0]; // @[LZD.scala 44:32]
  assign _T_1312 = _T_1311[3:2]; // @[LZD.scala 43:32]
  assign _T_1313 = _T_1312 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1314 = _T_1312[1]; // @[LZD.scala 39:21]
  assign _T_1315 = _T_1312[0]; // @[LZD.scala 39:30]
  assign _T_1316 = ~ _T_1315; // @[LZD.scala 39:27]
  assign _T_1317 = _T_1314 | _T_1316; // @[LZD.scala 39:25]
  assign _T_1318 = {_T_1313,_T_1317}; // @[Cat.scala 29:58]
  assign _T_1319 = _T_1311[1:0]; // @[LZD.scala 44:32]
  assign _T_1320 = _T_1319 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1321 = _T_1319[1]; // @[LZD.scala 39:21]
  assign _T_1322 = _T_1319[0]; // @[LZD.scala 39:30]
  assign _T_1323 = ~ _T_1322; // @[LZD.scala 39:27]
  assign _T_1324 = _T_1321 | _T_1323; // @[LZD.scala 39:25]
  assign _T_1325 = {_T_1320,_T_1324}; // @[Cat.scala 29:58]
  assign _T_1326 = _T_1318[1]; // @[Shift.scala 12:21]
  assign _T_1327 = _T_1325[1]; // @[Shift.scala 12:21]
  assign _T_1328 = _T_1326 | _T_1327; // @[LZD.scala 49:16]
  assign _T_1329 = ~ _T_1327; // @[LZD.scala 49:27]
  assign _T_1330 = _T_1326 | _T_1329; // @[LZD.scala 49:25]
  assign _T_1331 = _T_1318[0:0]; // @[LZD.scala 49:47]
  assign _T_1332 = _T_1325[0:0]; // @[LZD.scala 49:59]
  assign _T_1333 = _T_1326 ? _T_1331 : _T_1332; // @[LZD.scala 49:35]
  assign _T_1335 = {_T_1328,_T_1330,_T_1333}; // @[Cat.scala 29:58]
  assign _T_1336 = _T_1310[2]; // @[Shift.scala 12:21]
  assign _T_1337 = _T_1335[2]; // @[Shift.scala 12:21]
  assign _T_1338 = _T_1336 | _T_1337; // @[LZD.scala 49:16]
  assign _T_1339 = ~ _T_1337; // @[LZD.scala 49:27]
  assign _T_1340 = _T_1336 | _T_1339; // @[LZD.scala 49:25]
  assign _T_1341 = _T_1310[1:0]; // @[LZD.scala 49:47]
  assign _T_1342 = _T_1335[1:0]; // @[LZD.scala 49:59]
  assign _T_1343 = _T_1336 ? _T_1341 : _T_1342; // @[LZD.scala 49:35]
  assign _T_1345 = {_T_1338,_T_1340,_T_1343}; // @[Cat.scala 29:58]
  assign _T_1346 = _T_1284[7:0]; // @[LZD.scala 44:32]
  assign _T_1347 = _T_1346[7:4]; // @[LZD.scala 43:32]
  assign _T_1348 = _T_1347[3:2]; // @[LZD.scala 43:32]
  assign _T_1349 = _T_1348 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1350 = _T_1348[1]; // @[LZD.scala 39:21]
  assign _T_1351 = _T_1348[0]; // @[LZD.scala 39:30]
  assign _T_1352 = ~ _T_1351; // @[LZD.scala 39:27]
  assign _T_1353 = _T_1350 | _T_1352; // @[LZD.scala 39:25]
  assign _T_1354 = {_T_1349,_T_1353}; // @[Cat.scala 29:58]
  assign _T_1355 = _T_1347[1:0]; // @[LZD.scala 44:32]
  assign _T_1356 = _T_1355 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1357 = _T_1355[1]; // @[LZD.scala 39:21]
  assign _T_1358 = _T_1355[0]; // @[LZD.scala 39:30]
  assign _T_1359 = ~ _T_1358; // @[LZD.scala 39:27]
  assign _T_1360 = _T_1357 | _T_1359; // @[LZD.scala 39:25]
  assign _T_1361 = {_T_1356,_T_1360}; // @[Cat.scala 29:58]
  assign _T_1362 = _T_1354[1]; // @[Shift.scala 12:21]
  assign _T_1363 = _T_1361[1]; // @[Shift.scala 12:21]
  assign _T_1364 = _T_1362 | _T_1363; // @[LZD.scala 49:16]
  assign _T_1365 = ~ _T_1363; // @[LZD.scala 49:27]
  assign _T_1366 = _T_1362 | _T_1365; // @[LZD.scala 49:25]
  assign _T_1367 = _T_1354[0:0]; // @[LZD.scala 49:47]
  assign _T_1368 = _T_1361[0:0]; // @[LZD.scala 49:59]
  assign _T_1369 = _T_1362 ? _T_1367 : _T_1368; // @[LZD.scala 49:35]
  assign _T_1371 = {_T_1364,_T_1366,_T_1369}; // @[Cat.scala 29:58]
  assign _T_1372 = _T_1346[3:0]; // @[LZD.scala 44:32]
  assign _T_1373 = _T_1372[3:2]; // @[LZD.scala 43:32]
  assign _T_1374 = _T_1373 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1375 = _T_1373[1]; // @[LZD.scala 39:21]
  assign _T_1376 = _T_1373[0]; // @[LZD.scala 39:30]
  assign _T_1377 = ~ _T_1376; // @[LZD.scala 39:27]
  assign _T_1378 = _T_1375 | _T_1377; // @[LZD.scala 39:25]
  assign _T_1379 = {_T_1374,_T_1378}; // @[Cat.scala 29:58]
  assign _T_1380 = _T_1372[1:0]; // @[LZD.scala 44:32]
  assign _T_1381 = _T_1380 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1382 = _T_1380[1]; // @[LZD.scala 39:21]
  assign _T_1383 = _T_1380[0]; // @[LZD.scala 39:30]
  assign _T_1384 = ~ _T_1383; // @[LZD.scala 39:27]
  assign _T_1385 = _T_1382 | _T_1384; // @[LZD.scala 39:25]
  assign _T_1386 = {_T_1381,_T_1385}; // @[Cat.scala 29:58]
  assign _T_1387 = _T_1379[1]; // @[Shift.scala 12:21]
  assign _T_1388 = _T_1386[1]; // @[Shift.scala 12:21]
  assign _T_1389 = _T_1387 | _T_1388; // @[LZD.scala 49:16]
  assign _T_1390 = ~ _T_1388; // @[LZD.scala 49:27]
  assign _T_1391 = _T_1387 | _T_1390; // @[LZD.scala 49:25]
  assign _T_1392 = _T_1379[0:0]; // @[LZD.scala 49:47]
  assign _T_1393 = _T_1386[0:0]; // @[LZD.scala 49:59]
  assign _T_1394 = _T_1387 ? _T_1392 : _T_1393; // @[LZD.scala 49:35]
  assign _T_1396 = {_T_1389,_T_1391,_T_1394}; // @[Cat.scala 29:58]
  assign _T_1397 = _T_1371[2]; // @[Shift.scala 12:21]
  assign _T_1398 = _T_1396[2]; // @[Shift.scala 12:21]
  assign _T_1399 = _T_1397 | _T_1398; // @[LZD.scala 49:16]
  assign _T_1400 = ~ _T_1398; // @[LZD.scala 49:27]
  assign _T_1401 = _T_1397 | _T_1400; // @[LZD.scala 49:25]
  assign _T_1402 = _T_1371[1:0]; // @[LZD.scala 49:47]
  assign _T_1403 = _T_1396[1:0]; // @[LZD.scala 49:59]
  assign _T_1404 = _T_1397 ? _T_1402 : _T_1403; // @[LZD.scala 49:35]
  assign _T_1406 = {_T_1399,_T_1401,_T_1404}; // @[Cat.scala 29:58]
  assign _T_1407 = _T_1345[3]; // @[Shift.scala 12:21]
  assign _T_1408 = _T_1406[3]; // @[Shift.scala 12:21]
  assign _T_1409 = _T_1407 | _T_1408; // @[LZD.scala 49:16]
  assign _T_1410 = ~ _T_1408; // @[LZD.scala 49:27]
  assign _T_1411 = _T_1407 | _T_1410; // @[LZD.scala 49:25]
  assign _T_1412 = _T_1345[2:0]; // @[LZD.scala 49:47]
  assign _T_1413 = _T_1406[2:0]; // @[LZD.scala 49:59]
  assign _T_1414 = _T_1407 ? _T_1412 : _T_1413; // @[LZD.scala 49:35]
  assign _T_1416 = {_T_1409,_T_1411,_T_1414}; // @[Cat.scala 29:58]
  assign _T_1417 = _T_1283[0:0]; // @[LZD.scala 44:32]
  assign _T_1419 = _T_1416[4]; // @[Shift.scala 12:21]
  assign _T_1422 = {3'h7,_T_1417}; // @[Cat.scala 29:58]
  assign _T_1423 = _T_1416[3:0]; // @[LZD.scala 55:32]
  assign _T_1424 = _T_1419 ? _T_1423 : _T_1422; // @[LZD.scala 55:20]
  assign _T_1425 = {_T_1419,_T_1424}; // @[Cat.scala 29:58]
  assign _T_1426 = _T_1282[5]; // @[Shift.scala 12:21]
  assign _T_1428 = _T_1282[4:0]; // @[LZD.scala 55:32]
  assign _T_1429 = _T_1426 ? _T_1428 : _T_1425; // @[LZD.scala 55:20]
  assign sumLZD = {_T_1426,_T_1429}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 127:24]
  assign _T_1430 = signSumSig[47:0]; // @[PositFMA.scala 128:38]
  assign _T_1431 = shiftValue < 6'h30; // @[Shift.scala 16:24]
  assign _T_1433 = shiftValue[5]; // @[Shift.scala 12:21]
  assign _T_1434 = _T_1430[15:0]; // @[Shift.scala 64:52]
  assign _T_1436 = {_T_1434,32'h0}; // @[Cat.scala 29:58]
  assign _T_1437 = _T_1433 ? _T_1436 : _T_1430; // @[Shift.scala 64:27]
  assign _T_1438 = shiftValue[4:0]; // @[Shift.scala 66:70]
  assign _T_1439 = _T_1438[4]; // @[Shift.scala 12:21]
  assign _T_1440 = _T_1437[31:0]; // @[Shift.scala 64:52]
  assign _T_1442 = {_T_1440,16'h0}; // @[Cat.scala 29:58]
  assign _T_1443 = _T_1439 ? _T_1442 : _T_1437; // @[Shift.scala 64:27]
  assign _T_1444 = _T_1438[3:0]; // @[Shift.scala 66:70]
  assign _T_1445 = _T_1444[3]; // @[Shift.scala 12:21]
  assign _T_1446 = _T_1443[39:0]; // @[Shift.scala 64:52]
  assign _T_1448 = {_T_1446,8'h0}; // @[Cat.scala 29:58]
  assign _T_1449 = _T_1445 ? _T_1448 : _T_1443; // @[Shift.scala 64:27]
  assign _T_1450 = _T_1444[2:0]; // @[Shift.scala 66:70]
  assign _T_1451 = _T_1450[2]; // @[Shift.scala 12:21]
  assign _T_1452 = _T_1449[43:0]; // @[Shift.scala 64:52]
  assign _T_1454 = {_T_1452,4'h0}; // @[Cat.scala 29:58]
  assign _T_1455 = _T_1451 ? _T_1454 : _T_1449; // @[Shift.scala 64:27]
  assign _T_1456 = _T_1450[1:0]; // @[Shift.scala 66:70]
  assign _T_1457 = _T_1456[1]; // @[Shift.scala 12:21]
  assign _T_1458 = _T_1455[45:0]; // @[Shift.scala 64:52]
  assign _T_1460 = {_T_1458,2'h0}; // @[Cat.scala 29:58]
  assign _T_1461 = _T_1457 ? _T_1460 : _T_1455; // @[Shift.scala 64:27]
  assign _T_1462 = _T_1456[0:0]; // @[Shift.scala 66:70]
  assign _T_1464 = _T_1461[46:0]; // @[Shift.scala 64:52]
  assign _T_1465 = {_T_1464,1'h0}; // @[Cat.scala 29:58]
  assign _T_1466 = _T_1462 ? _T_1465 : _T_1461; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_1431 ? _T_1466 : 48'h0; // @[Shift.scala 16:10]
  assign _T_1468 = $signed(greaterScale) + $signed(10'sh2); // @[PositFMA.scala 131:36]
  assign _T_1469 = $signed(_T_1468); // @[PositFMA.scala 131:36]
  assign _T_1470 = {1'h1,_T_1426,_T_1429}; // @[Cat.scala 29:58]
  assign _T_1471 = $signed(_T_1470); // @[PositFMA.scala 131:61]
  assign _GEN_20 = {{3{_T_1471[6]}},_T_1471}; // @[PositFMA.scala 131:42]
  assign _T_1473 = $signed(_T_1469) + $signed(_GEN_20); // @[PositFMA.scala 131:42]
  assign sumScale = $signed(_T_1473); // @[PositFMA.scala 131:42]
  assign sumFrac = normalFracTmp[47:25]; // @[PositFMA.scala 132:41]
  assign grsTmp = normalFracTmp[24:0]; // @[PositFMA.scala 135:41]
  assign _T_1474 = grsTmp[24:23]; // @[PositFMA.scala 138:40]
  assign _T_1475 = grsTmp[22:0]; // @[PositFMA.scala 138:56]
  assign _T_1476 = _T_1475 != 23'h0; // @[PositFMA.scala 138:60]
  assign underflow = $signed(sumScale) < $signed(-10'shd8); // @[PositFMA.scala 145:32]
  assign overflow = $signed(sumScale) > $signed(10'shd8); // @[PositFMA.scala 146:32]
  assign _T_1477 = signSumSig != 50'h0; // @[PositFMA.scala 155:32]
  assign decF_isZero = ~ _T_1477; // @[PositFMA.scala 155:20]
  assign _T_1479 = underflow ? $signed(-10'shd8) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_1480 = overflow ? $signed(10'shd8) : $signed(_T_1479); // @[Mux.scala 87:16]
  assign _GEN_21 = _T_1480[8:0]; // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  assign decF_scale = $signed(_GEN_21); // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  assign _T_1481 = decF_scale[2:0]; // @[convert.scala 46:61]
  assign _T_1482 = ~ _T_1481; // @[convert.scala 46:52]
  assign _T_1484 = sumSign ? _T_1482 : _T_1481; // @[convert.scala 46:42]
  assign _T_1485 = decF_scale[8:3]; // @[convert.scala 48:34]
  assign _T_1486 = _T_1485[5:5]; // @[convert.scala 49:36]
  assign _T_1488 = ~ _T_1485; // @[convert.scala 50:36]
  assign _T_1489 = $signed(_T_1488); // @[convert.scala 50:36]
  assign _T_1490 = _T_1486 ? $signed(_T_1489) : $signed(_T_1485); // @[convert.scala 50:28]
  assign _T_1491 = _T_1486 ^ sumSign; // @[convert.scala 51:31]
  assign _T_1492 = ~ _T_1491; // @[convert.scala 52:43]
  assign _T_1496 = {_T_1492,_T_1491,_T_1484,sumFrac,_T_1474,_T_1476}; // @[Cat.scala 29:58]
  assign _T_1497 = $unsigned(_T_1490); // @[Shift.scala 39:17]
  assign _T_1498 = _T_1497 < 6'h1f; // @[Shift.scala 39:24]
  assign _T_1499 = _T_1490[4:0]; // @[Shift.scala 40:44]
  assign _T_1500 = _T_1496[30:16]; // @[Shift.scala 90:30]
  assign _T_1501 = _T_1496[15:0]; // @[Shift.scala 90:48]
  assign _T_1502 = _T_1501 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{14'd0}, _T_1502}; // @[Shift.scala 90:39]
  assign _T_1503 = _T_1500 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_1504 = _T_1499[4]; // @[Shift.scala 12:21]
  assign _T_1505 = _T_1496[30]; // @[Shift.scala 12:21]
  assign _T_1507 = _T_1505 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_1508 = {_T_1507,_T_1503}; // @[Cat.scala 29:58]
  assign _T_1509 = _T_1504 ? _T_1508 : _T_1496; // @[Shift.scala 91:22]
  assign _T_1510 = _T_1499[3:0]; // @[Shift.scala 92:77]
  assign _T_1511 = _T_1509[30:8]; // @[Shift.scala 90:30]
  assign _T_1512 = _T_1509[7:0]; // @[Shift.scala 90:48]
  assign _T_1513 = _T_1512 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{22'd0}, _T_1513}; // @[Shift.scala 90:39]
  assign _T_1514 = _T_1511 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_1515 = _T_1510[3]; // @[Shift.scala 12:21]
  assign _T_1516 = _T_1509[30]; // @[Shift.scala 12:21]
  assign _T_1518 = _T_1516 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_1519 = {_T_1518,_T_1514}; // @[Cat.scala 29:58]
  assign _T_1520 = _T_1515 ? _T_1519 : _T_1509; // @[Shift.scala 91:22]
  assign _T_1521 = _T_1510[2:0]; // @[Shift.scala 92:77]
  assign _T_1522 = _T_1520[30:4]; // @[Shift.scala 90:30]
  assign _T_1523 = _T_1520[3:0]; // @[Shift.scala 90:48]
  assign _T_1524 = _T_1523 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_24 = {{26'd0}, _T_1524}; // @[Shift.scala 90:39]
  assign _T_1525 = _T_1522 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_1526 = _T_1521[2]; // @[Shift.scala 12:21]
  assign _T_1527 = _T_1520[30]; // @[Shift.scala 12:21]
  assign _T_1529 = _T_1527 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_1530 = {_T_1529,_T_1525}; // @[Cat.scala 29:58]
  assign _T_1531 = _T_1526 ? _T_1530 : _T_1520; // @[Shift.scala 91:22]
  assign _T_1532 = _T_1521[1:0]; // @[Shift.scala 92:77]
  assign _T_1533 = _T_1531[30:2]; // @[Shift.scala 90:30]
  assign _T_1534 = _T_1531[1:0]; // @[Shift.scala 90:48]
  assign _T_1535 = _T_1534 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_25 = {{28'd0}, _T_1535}; // @[Shift.scala 90:39]
  assign _T_1536 = _T_1533 | _GEN_25; // @[Shift.scala 90:39]
  assign _T_1537 = _T_1532[1]; // @[Shift.scala 12:21]
  assign _T_1538 = _T_1531[30]; // @[Shift.scala 12:21]
  assign _T_1540 = _T_1538 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_1541 = {_T_1540,_T_1536}; // @[Cat.scala 29:58]
  assign _T_1542 = _T_1537 ? _T_1541 : _T_1531; // @[Shift.scala 91:22]
  assign _T_1543 = _T_1532[0:0]; // @[Shift.scala 92:77]
  assign _T_1544 = _T_1542[30:1]; // @[Shift.scala 90:30]
  assign _T_1545 = _T_1542[0:0]; // @[Shift.scala 90:48]
  assign _GEN_26 = {{29'd0}, _T_1545}; // @[Shift.scala 90:39]
  assign _T_1547 = _T_1544 | _GEN_26; // @[Shift.scala 90:39]
  assign _T_1549 = _T_1542[30]; // @[Shift.scala 12:21]
  assign _T_1550 = {_T_1549,_T_1547}; // @[Cat.scala 29:58]
  assign _T_1551 = _T_1543 ? _T_1550 : _T_1542; // @[Shift.scala 91:22]
  assign _T_1554 = _T_1505 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 71:12]
  assign _T_1555 = _T_1498 ? _T_1551 : _T_1554; // @[Shift.scala 39:10]
  assign _T_1556 = _T_1555[3]; // @[convert.scala 55:31]
  assign _T_1557 = _T_1555[2]; // @[convert.scala 56:31]
  assign _T_1558 = _T_1555[1]; // @[convert.scala 57:31]
  assign _T_1559 = _T_1555[0]; // @[convert.scala 58:31]
  assign _T_1560 = _T_1555[30:3]; // @[convert.scala 59:69]
  assign _T_1561 = _T_1560 != 28'h0; // @[convert.scala 59:81]
  assign _T_1562 = ~ _T_1561; // @[convert.scala 59:50]
  assign _T_1564 = _T_1560 == 28'hfffffff; // @[convert.scala 60:81]
  assign _T_1565 = _T_1556 | _T_1558; // @[convert.scala 61:44]
  assign _T_1566 = _T_1565 | _T_1559; // @[convert.scala 61:52]
  assign _T_1567 = _T_1557 & _T_1566; // @[convert.scala 61:36]
  assign _T_1568 = ~ _T_1564; // @[convert.scala 62:63]
  assign _T_1569 = _T_1568 & _T_1567; // @[convert.scala 62:103]
  assign _T_1570 = _T_1562 | _T_1569; // @[convert.scala 62:60]
  assign _GEN_27 = {{27'd0}, _T_1570}; // @[convert.scala 63:56]
  assign _T_1573 = _T_1560 + _GEN_27; // @[convert.scala 63:56]
  assign _T_1574 = {sumSign,_T_1573}; // @[Cat.scala 29:58]
  assign io_F = _T_1582; // @[PositFMA.scala 175:15]
  assign io_outValid = _T_1578; // @[PositFMA.scala 174:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  mulSig_phase2 = _RAND_1[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[22:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1578 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1582 = _RAND_9[28:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_583;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_1578 <= 1'h0;
    end else begin
      _T_1578 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_1582 <= 29'h10000000;
      end else begin
        if (decF_isZero) begin
          _T_1582 <= 29'h0;
        end else begin
          _T_1582 <= _T_1574;
        end
      end
    end
  end
endmodule
