module PositDivSqrter30_3(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [29:0] io_A,
  input  [29:0] io_B,
  output        io_diviValid,
  output        io_sqrtValid,
  output        io_invalidExc,
  output [29:0] io_Q
);
  reg [4:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [9:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [23:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [27:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [27:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [27:0] _T_4; // @[convert.scala 19:24]
  wire [27:0] _T_5; // @[convert.scala 19:43]
  wire [27:0] _T_6; // @[convert.scala 19:39]
  wire [15:0] _T_7; // @[LZD.scala 43:32]
  wire [7:0] _T_8; // @[LZD.scala 43:32]
  wire [3:0] _T_9; // @[LZD.scala 43:32]
  wire [1:0] _T_10; // @[LZD.scala 43:32]
  wire  _T_11; // @[LZD.scala 39:14]
  wire  _T_12; // @[LZD.scala 39:21]
  wire  _T_13; // @[LZD.scala 39:30]
  wire  _T_14; // @[LZD.scala 39:27]
  wire  _T_15; // @[LZD.scala 39:25]
  wire [1:0] _T_16; // @[Cat.scala 29:58]
  wire [1:0] _T_17; // @[LZD.scala 44:32]
  wire  _T_18; // @[LZD.scala 39:14]
  wire  _T_19; // @[LZD.scala 39:21]
  wire  _T_20; // @[LZD.scala 39:30]
  wire  _T_21; // @[LZD.scala 39:27]
  wire  _T_22; // @[LZD.scala 39:25]
  wire [1:0] _T_23; // @[Cat.scala 29:58]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[Shift.scala 12:21]
  wire  _T_26; // @[LZD.scala 49:16]
  wire  _T_27; // @[LZD.scala 49:27]
  wire  _T_28; // @[LZD.scala 49:25]
  wire  _T_29; // @[LZD.scala 49:47]
  wire  _T_30; // @[LZD.scala 49:59]
  wire  _T_31; // @[LZD.scala 49:35]
  wire [2:0] _T_33; // @[Cat.scala 29:58]
  wire [3:0] _T_34; // @[LZD.scala 44:32]
  wire [1:0] _T_35; // @[LZD.scala 43:32]
  wire  _T_36; // @[LZD.scala 39:14]
  wire  _T_37; // @[LZD.scala 39:21]
  wire  _T_38; // @[LZD.scala 39:30]
  wire  _T_39; // @[LZD.scala 39:27]
  wire  _T_40; // @[LZD.scala 39:25]
  wire [1:0] _T_41; // @[Cat.scala 29:58]
  wire [1:0] _T_42; // @[LZD.scala 44:32]
  wire  _T_43; // @[LZD.scala 39:14]
  wire  _T_44; // @[LZD.scala 39:21]
  wire  _T_45; // @[LZD.scala 39:30]
  wire  _T_46; // @[LZD.scala 39:27]
  wire  _T_47; // @[LZD.scala 39:25]
  wire [1:0] _T_48; // @[Cat.scala 29:58]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[Shift.scala 12:21]
  wire  _T_51; // @[LZD.scala 49:16]
  wire  _T_52; // @[LZD.scala 49:27]
  wire  _T_53; // @[LZD.scala 49:25]
  wire  _T_54; // @[LZD.scala 49:47]
  wire  _T_55; // @[LZD.scala 49:59]
  wire  _T_56; // @[LZD.scala 49:35]
  wire [2:0] _T_58; // @[Cat.scala 29:58]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[LZD.scala 49:16]
  wire  _T_62; // @[LZD.scala 49:27]
  wire  _T_63; // @[LZD.scala 49:25]
  wire [1:0] _T_64; // @[LZD.scala 49:47]
  wire [1:0] _T_65; // @[LZD.scala 49:59]
  wire [1:0] _T_66; // @[LZD.scala 49:35]
  wire [3:0] _T_68; // @[Cat.scala 29:58]
  wire [7:0] _T_69; // @[LZD.scala 44:32]
  wire [3:0] _T_70; // @[LZD.scala 43:32]
  wire [1:0] _T_71; // @[LZD.scala 43:32]
  wire  _T_72; // @[LZD.scala 39:14]
  wire  _T_73; // @[LZD.scala 39:21]
  wire  _T_74; // @[LZD.scala 39:30]
  wire  _T_75; // @[LZD.scala 39:27]
  wire  _T_76; // @[LZD.scala 39:25]
  wire [1:0] _T_77; // @[Cat.scala 29:58]
  wire [1:0] _T_78; // @[LZD.scala 44:32]
  wire  _T_79; // @[LZD.scala 39:14]
  wire  _T_80; // @[LZD.scala 39:21]
  wire  _T_81; // @[LZD.scala 39:30]
  wire  _T_82; // @[LZD.scala 39:27]
  wire  _T_83; // @[LZD.scala 39:25]
  wire [1:0] _T_84; // @[Cat.scala 29:58]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[Shift.scala 12:21]
  wire  _T_87; // @[LZD.scala 49:16]
  wire  _T_88; // @[LZD.scala 49:27]
  wire  _T_89; // @[LZD.scala 49:25]
  wire  _T_90; // @[LZD.scala 49:47]
  wire  _T_91; // @[LZD.scala 49:59]
  wire  _T_92; // @[LZD.scala 49:35]
  wire [2:0] _T_94; // @[Cat.scala 29:58]
  wire [3:0] _T_95; // @[LZD.scala 44:32]
  wire [1:0] _T_96; // @[LZD.scala 43:32]
  wire  _T_97; // @[LZD.scala 39:14]
  wire  _T_98; // @[LZD.scala 39:21]
  wire  _T_99; // @[LZD.scala 39:30]
  wire  _T_100; // @[LZD.scala 39:27]
  wire  _T_101; // @[LZD.scala 39:25]
  wire [1:0] _T_102; // @[Cat.scala 29:58]
  wire [1:0] _T_103; // @[LZD.scala 44:32]
  wire  _T_104; // @[LZD.scala 39:14]
  wire  _T_105; // @[LZD.scala 39:21]
  wire  _T_106; // @[LZD.scala 39:30]
  wire  _T_107; // @[LZD.scala 39:27]
  wire  _T_108; // @[LZD.scala 39:25]
  wire [1:0] _T_109; // @[Cat.scala 29:58]
  wire  _T_110; // @[Shift.scala 12:21]
  wire  _T_111; // @[Shift.scala 12:21]
  wire  _T_112; // @[LZD.scala 49:16]
  wire  _T_113; // @[LZD.scala 49:27]
  wire  _T_114; // @[LZD.scala 49:25]
  wire  _T_115; // @[LZD.scala 49:47]
  wire  _T_116; // @[LZD.scala 49:59]
  wire  _T_117; // @[LZD.scala 49:35]
  wire [2:0] _T_119; // @[Cat.scala 29:58]
  wire  _T_120; // @[Shift.scala 12:21]
  wire  _T_121; // @[Shift.scala 12:21]
  wire  _T_122; // @[LZD.scala 49:16]
  wire  _T_123; // @[LZD.scala 49:27]
  wire  _T_124; // @[LZD.scala 49:25]
  wire [1:0] _T_125; // @[LZD.scala 49:47]
  wire [1:0] _T_126; // @[LZD.scala 49:59]
  wire [1:0] _T_127; // @[LZD.scala 49:35]
  wire [3:0] _T_129; // @[Cat.scala 29:58]
  wire  _T_130; // @[Shift.scala 12:21]
  wire  _T_131; // @[Shift.scala 12:21]
  wire  _T_132; // @[LZD.scala 49:16]
  wire  _T_133; // @[LZD.scala 49:27]
  wire  _T_134; // @[LZD.scala 49:25]
  wire [2:0] _T_135; // @[LZD.scala 49:47]
  wire [2:0] _T_136; // @[LZD.scala 49:59]
  wire [2:0] _T_137; // @[LZD.scala 49:35]
  wire [4:0] _T_139; // @[Cat.scala 29:58]
  wire [11:0] _T_140; // @[LZD.scala 44:32]
  wire [7:0] _T_141; // @[LZD.scala 43:32]
  wire [3:0] _T_142; // @[LZD.scala 43:32]
  wire [1:0] _T_143; // @[LZD.scala 43:32]
  wire  _T_144; // @[LZD.scala 39:14]
  wire  _T_145; // @[LZD.scala 39:21]
  wire  _T_146; // @[LZD.scala 39:30]
  wire  _T_147; // @[LZD.scala 39:27]
  wire  _T_148; // @[LZD.scala 39:25]
  wire [1:0] _T_149; // @[Cat.scala 29:58]
  wire [1:0] _T_150; // @[LZD.scala 44:32]
  wire  _T_151; // @[LZD.scala 39:14]
  wire  _T_152; // @[LZD.scala 39:21]
  wire  _T_153; // @[LZD.scala 39:30]
  wire  _T_154; // @[LZD.scala 39:27]
  wire  _T_155; // @[LZD.scala 39:25]
  wire [1:0] _T_156; // @[Cat.scala 29:58]
  wire  _T_157; // @[Shift.scala 12:21]
  wire  _T_158; // @[Shift.scala 12:21]
  wire  _T_159; // @[LZD.scala 49:16]
  wire  _T_160; // @[LZD.scala 49:27]
  wire  _T_161; // @[LZD.scala 49:25]
  wire  _T_162; // @[LZD.scala 49:47]
  wire  _T_163; // @[LZD.scala 49:59]
  wire  _T_164; // @[LZD.scala 49:35]
  wire [2:0] _T_166; // @[Cat.scala 29:58]
  wire [3:0] _T_167; // @[LZD.scala 44:32]
  wire [1:0] _T_168; // @[LZD.scala 43:32]
  wire  _T_169; // @[LZD.scala 39:14]
  wire  _T_170; // @[LZD.scala 39:21]
  wire  _T_171; // @[LZD.scala 39:30]
  wire  _T_172; // @[LZD.scala 39:27]
  wire  _T_173; // @[LZD.scala 39:25]
  wire [1:0] _T_174; // @[Cat.scala 29:58]
  wire [1:0] _T_175; // @[LZD.scala 44:32]
  wire  _T_176; // @[LZD.scala 39:14]
  wire  _T_177; // @[LZD.scala 39:21]
  wire  _T_178; // @[LZD.scala 39:30]
  wire  _T_179; // @[LZD.scala 39:27]
  wire  _T_180; // @[LZD.scala 39:25]
  wire [1:0] _T_181; // @[Cat.scala 29:58]
  wire  _T_182; // @[Shift.scala 12:21]
  wire  _T_183; // @[Shift.scala 12:21]
  wire  _T_184; // @[LZD.scala 49:16]
  wire  _T_185; // @[LZD.scala 49:27]
  wire  _T_186; // @[LZD.scala 49:25]
  wire  _T_187; // @[LZD.scala 49:47]
  wire  _T_188; // @[LZD.scala 49:59]
  wire  _T_189; // @[LZD.scala 49:35]
  wire [2:0] _T_191; // @[Cat.scala 29:58]
  wire  _T_192; // @[Shift.scala 12:21]
  wire  _T_193; // @[Shift.scala 12:21]
  wire  _T_194; // @[LZD.scala 49:16]
  wire  _T_195; // @[LZD.scala 49:27]
  wire  _T_196; // @[LZD.scala 49:25]
  wire [1:0] _T_197; // @[LZD.scala 49:47]
  wire [1:0] _T_198; // @[LZD.scala 49:59]
  wire [1:0] _T_199; // @[LZD.scala 49:35]
  wire [3:0] _T_201; // @[Cat.scala 29:58]
  wire [3:0] _T_202; // @[LZD.scala 44:32]
  wire [1:0] _T_203; // @[LZD.scala 43:32]
  wire  _T_204; // @[LZD.scala 39:14]
  wire  _T_205; // @[LZD.scala 39:21]
  wire  _T_206; // @[LZD.scala 39:30]
  wire  _T_207; // @[LZD.scala 39:27]
  wire  _T_208; // @[LZD.scala 39:25]
  wire [1:0] _T_209; // @[Cat.scala 29:58]
  wire [1:0] _T_210; // @[LZD.scala 44:32]
  wire  _T_211; // @[LZD.scala 39:14]
  wire  _T_212; // @[LZD.scala 39:21]
  wire  _T_213; // @[LZD.scala 39:30]
  wire  _T_214; // @[LZD.scala 39:27]
  wire  _T_215; // @[LZD.scala 39:25]
  wire [1:0] _T_216; // @[Cat.scala 29:58]
  wire  _T_217; // @[Shift.scala 12:21]
  wire  _T_218; // @[Shift.scala 12:21]
  wire  _T_219; // @[LZD.scala 49:16]
  wire  _T_220; // @[LZD.scala 49:27]
  wire  _T_221; // @[LZD.scala 49:25]
  wire  _T_222; // @[LZD.scala 49:47]
  wire  _T_223; // @[LZD.scala 49:59]
  wire  _T_224; // @[LZD.scala 49:35]
  wire [2:0] _T_226; // @[Cat.scala 29:58]
  wire  _T_227; // @[Shift.scala 12:21]
  wire [2:0] _T_229; // @[LZD.scala 55:32]
  wire [2:0] _T_230; // @[LZD.scala 55:20]
  wire [3:0] _T_231; // @[Cat.scala 29:58]
  wire  _T_232; // @[Shift.scala 12:21]
  wire [3:0] _T_234; // @[LZD.scala 55:32]
  wire [3:0] _T_235; // @[LZD.scala 55:20]
  wire [4:0] _T_236; // @[Cat.scala 29:58]
  wire [4:0] _T_237; // @[convert.scala 21:22]
  wire [26:0] _T_238; // @[convert.scala 22:36]
  wire  _T_239; // @[Shift.scala 16:24]
  wire  _T_241; // @[Shift.scala 12:21]
  wire [10:0] _T_242; // @[Shift.scala 64:52]
  wire [26:0] _T_244; // @[Cat.scala 29:58]
  wire [26:0] _T_245; // @[Shift.scala 64:27]
  wire [3:0] _T_246; // @[Shift.scala 66:70]
  wire  _T_247; // @[Shift.scala 12:21]
  wire [18:0] _T_248; // @[Shift.scala 64:52]
  wire [26:0] _T_250; // @[Cat.scala 29:58]
  wire [26:0] _T_251; // @[Shift.scala 64:27]
  wire [2:0] _T_252; // @[Shift.scala 66:70]
  wire  _T_253; // @[Shift.scala 12:21]
  wire [22:0] _T_254; // @[Shift.scala 64:52]
  wire [26:0] _T_256; // @[Cat.scala 29:58]
  wire [26:0] _T_257; // @[Shift.scala 64:27]
  wire [1:0] _T_258; // @[Shift.scala 66:70]
  wire  _T_259; // @[Shift.scala 12:21]
  wire [24:0] _T_260; // @[Shift.scala 64:52]
  wire [26:0] _T_262; // @[Cat.scala 29:58]
  wire [26:0] _T_263; // @[Shift.scala 64:27]
  wire  _T_264; // @[Shift.scala 66:70]
  wire [25:0] _T_266; // @[Shift.scala 64:52]
  wire [26:0] _T_267; // @[Cat.scala 29:58]
  wire [26:0] _T_268; // @[Shift.scala 64:27]
  wire [26:0] _T_269; // @[Shift.scala 16:10]
  wire [2:0] _T_270; // @[convert.scala 23:34]
  wire [23:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_272; // @[convert.scala 25:26]
  wire [4:0] _T_274; // @[convert.scala 25:42]
  wire [2:0] _T_277; // @[convert.scala 26:67]
  wire [2:0] _T_278; // @[convert.scala 26:51]
  wire [8:0] _T_279; // @[Cat.scala 29:58]
  wire [28:0] _T_281; // @[convert.scala 29:56]
  wire  _T_282; // @[convert.scala 29:60]
  wire  _T_283; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_286; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [8:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_295; // @[convert.scala 18:24]
  wire  _T_296; // @[convert.scala 18:40]
  wire  _T_297; // @[convert.scala 18:36]
  wire [27:0] _T_298; // @[convert.scala 19:24]
  wire [27:0] _T_299; // @[convert.scala 19:43]
  wire [27:0] _T_300; // @[convert.scala 19:39]
  wire [15:0] _T_301; // @[LZD.scala 43:32]
  wire [7:0] _T_302; // @[LZD.scala 43:32]
  wire [3:0] _T_303; // @[LZD.scala 43:32]
  wire [1:0] _T_304; // @[LZD.scala 43:32]
  wire  _T_305; // @[LZD.scala 39:14]
  wire  _T_306; // @[LZD.scala 39:21]
  wire  _T_307; // @[LZD.scala 39:30]
  wire  _T_308; // @[LZD.scala 39:27]
  wire  _T_309; // @[LZD.scala 39:25]
  wire [1:0] _T_310; // @[Cat.scala 29:58]
  wire [1:0] _T_311; // @[LZD.scala 44:32]
  wire  _T_312; // @[LZD.scala 39:14]
  wire  _T_313; // @[LZD.scala 39:21]
  wire  _T_314; // @[LZD.scala 39:30]
  wire  _T_315; // @[LZD.scala 39:27]
  wire  _T_316; // @[LZD.scala 39:25]
  wire [1:0] _T_317; // @[Cat.scala 29:58]
  wire  _T_318; // @[Shift.scala 12:21]
  wire  _T_319; // @[Shift.scala 12:21]
  wire  _T_320; // @[LZD.scala 49:16]
  wire  _T_321; // @[LZD.scala 49:27]
  wire  _T_322; // @[LZD.scala 49:25]
  wire  _T_323; // @[LZD.scala 49:47]
  wire  _T_324; // @[LZD.scala 49:59]
  wire  _T_325; // @[LZD.scala 49:35]
  wire [2:0] _T_327; // @[Cat.scala 29:58]
  wire [3:0] _T_328; // @[LZD.scala 44:32]
  wire [1:0] _T_329; // @[LZD.scala 43:32]
  wire  _T_330; // @[LZD.scala 39:14]
  wire  _T_331; // @[LZD.scala 39:21]
  wire  _T_332; // @[LZD.scala 39:30]
  wire  _T_333; // @[LZD.scala 39:27]
  wire  _T_334; // @[LZD.scala 39:25]
  wire [1:0] _T_335; // @[Cat.scala 29:58]
  wire [1:0] _T_336; // @[LZD.scala 44:32]
  wire  _T_337; // @[LZD.scala 39:14]
  wire  _T_338; // @[LZD.scala 39:21]
  wire  _T_339; // @[LZD.scala 39:30]
  wire  _T_340; // @[LZD.scala 39:27]
  wire  _T_341; // @[LZD.scala 39:25]
  wire [1:0] _T_342; // @[Cat.scala 29:58]
  wire  _T_343; // @[Shift.scala 12:21]
  wire  _T_344; // @[Shift.scala 12:21]
  wire  _T_345; // @[LZD.scala 49:16]
  wire  _T_346; // @[LZD.scala 49:27]
  wire  _T_347; // @[LZD.scala 49:25]
  wire  _T_348; // @[LZD.scala 49:47]
  wire  _T_349; // @[LZD.scala 49:59]
  wire  _T_350; // @[LZD.scala 49:35]
  wire [2:0] _T_352; // @[Cat.scala 29:58]
  wire  _T_353; // @[Shift.scala 12:21]
  wire  _T_354; // @[Shift.scala 12:21]
  wire  _T_355; // @[LZD.scala 49:16]
  wire  _T_356; // @[LZD.scala 49:27]
  wire  _T_357; // @[LZD.scala 49:25]
  wire [1:0] _T_358; // @[LZD.scala 49:47]
  wire [1:0] _T_359; // @[LZD.scala 49:59]
  wire [1:0] _T_360; // @[LZD.scala 49:35]
  wire [3:0] _T_362; // @[Cat.scala 29:58]
  wire [7:0] _T_363; // @[LZD.scala 44:32]
  wire [3:0] _T_364; // @[LZD.scala 43:32]
  wire [1:0] _T_365; // @[LZD.scala 43:32]
  wire  _T_366; // @[LZD.scala 39:14]
  wire  _T_367; // @[LZD.scala 39:21]
  wire  _T_368; // @[LZD.scala 39:30]
  wire  _T_369; // @[LZD.scala 39:27]
  wire  _T_370; // @[LZD.scala 39:25]
  wire [1:0] _T_371; // @[Cat.scala 29:58]
  wire [1:0] _T_372; // @[LZD.scala 44:32]
  wire  _T_373; // @[LZD.scala 39:14]
  wire  _T_374; // @[LZD.scala 39:21]
  wire  _T_375; // @[LZD.scala 39:30]
  wire  _T_376; // @[LZD.scala 39:27]
  wire  _T_377; // @[LZD.scala 39:25]
  wire [1:0] _T_378; // @[Cat.scala 29:58]
  wire  _T_379; // @[Shift.scala 12:21]
  wire  _T_380; // @[Shift.scala 12:21]
  wire  _T_381; // @[LZD.scala 49:16]
  wire  _T_382; // @[LZD.scala 49:27]
  wire  _T_383; // @[LZD.scala 49:25]
  wire  _T_384; // @[LZD.scala 49:47]
  wire  _T_385; // @[LZD.scala 49:59]
  wire  _T_386; // @[LZD.scala 49:35]
  wire [2:0] _T_388; // @[Cat.scala 29:58]
  wire [3:0] _T_389; // @[LZD.scala 44:32]
  wire [1:0] _T_390; // @[LZD.scala 43:32]
  wire  _T_391; // @[LZD.scala 39:14]
  wire  _T_392; // @[LZD.scala 39:21]
  wire  _T_393; // @[LZD.scala 39:30]
  wire  _T_394; // @[LZD.scala 39:27]
  wire  _T_395; // @[LZD.scala 39:25]
  wire [1:0] _T_396; // @[Cat.scala 29:58]
  wire [1:0] _T_397; // @[LZD.scala 44:32]
  wire  _T_398; // @[LZD.scala 39:14]
  wire  _T_399; // @[LZD.scala 39:21]
  wire  _T_400; // @[LZD.scala 39:30]
  wire  _T_401; // @[LZD.scala 39:27]
  wire  _T_402; // @[LZD.scala 39:25]
  wire [1:0] _T_403; // @[Cat.scala 29:58]
  wire  _T_404; // @[Shift.scala 12:21]
  wire  _T_405; // @[Shift.scala 12:21]
  wire  _T_406; // @[LZD.scala 49:16]
  wire  _T_407; // @[LZD.scala 49:27]
  wire  _T_408; // @[LZD.scala 49:25]
  wire  _T_409; // @[LZD.scala 49:47]
  wire  _T_410; // @[LZD.scala 49:59]
  wire  _T_411; // @[LZD.scala 49:35]
  wire [2:0] _T_413; // @[Cat.scala 29:58]
  wire  _T_414; // @[Shift.scala 12:21]
  wire  _T_415; // @[Shift.scala 12:21]
  wire  _T_416; // @[LZD.scala 49:16]
  wire  _T_417; // @[LZD.scala 49:27]
  wire  _T_418; // @[LZD.scala 49:25]
  wire [1:0] _T_419; // @[LZD.scala 49:47]
  wire [1:0] _T_420; // @[LZD.scala 49:59]
  wire [1:0] _T_421; // @[LZD.scala 49:35]
  wire [3:0] _T_423; // @[Cat.scala 29:58]
  wire  _T_424; // @[Shift.scala 12:21]
  wire  _T_425; // @[Shift.scala 12:21]
  wire  _T_426; // @[LZD.scala 49:16]
  wire  _T_427; // @[LZD.scala 49:27]
  wire  _T_428; // @[LZD.scala 49:25]
  wire [2:0] _T_429; // @[LZD.scala 49:47]
  wire [2:0] _T_430; // @[LZD.scala 49:59]
  wire [2:0] _T_431; // @[LZD.scala 49:35]
  wire [4:0] _T_433; // @[Cat.scala 29:58]
  wire [11:0] _T_434; // @[LZD.scala 44:32]
  wire [7:0] _T_435; // @[LZD.scala 43:32]
  wire [3:0] _T_436; // @[LZD.scala 43:32]
  wire [1:0] _T_437; // @[LZD.scala 43:32]
  wire  _T_438; // @[LZD.scala 39:14]
  wire  _T_439; // @[LZD.scala 39:21]
  wire  _T_440; // @[LZD.scala 39:30]
  wire  _T_441; // @[LZD.scala 39:27]
  wire  _T_442; // @[LZD.scala 39:25]
  wire [1:0] _T_443; // @[Cat.scala 29:58]
  wire [1:0] _T_444; // @[LZD.scala 44:32]
  wire  _T_445; // @[LZD.scala 39:14]
  wire  _T_446; // @[LZD.scala 39:21]
  wire  _T_447; // @[LZD.scala 39:30]
  wire  _T_448; // @[LZD.scala 39:27]
  wire  _T_449; // @[LZD.scala 39:25]
  wire [1:0] _T_450; // @[Cat.scala 29:58]
  wire  _T_451; // @[Shift.scala 12:21]
  wire  _T_452; // @[Shift.scala 12:21]
  wire  _T_453; // @[LZD.scala 49:16]
  wire  _T_454; // @[LZD.scala 49:27]
  wire  _T_455; // @[LZD.scala 49:25]
  wire  _T_456; // @[LZD.scala 49:47]
  wire  _T_457; // @[LZD.scala 49:59]
  wire  _T_458; // @[LZD.scala 49:35]
  wire [2:0] _T_460; // @[Cat.scala 29:58]
  wire [3:0] _T_461; // @[LZD.scala 44:32]
  wire [1:0] _T_462; // @[LZD.scala 43:32]
  wire  _T_463; // @[LZD.scala 39:14]
  wire  _T_464; // @[LZD.scala 39:21]
  wire  _T_465; // @[LZD.scala 39:30]
  wire  _T_466; // @[LZD.scala 39:27]
  wire  _T_467; // @[LZD.scala 39:25]
  wire [1:0] _T_468; // @[Cat.scala 29:58]
  wire [1:0] _T_469; // @[LZD.scala 44:32]
  wire  _T_470; // @[LZD.scala 39:14]
  wire  _T_471; // @[LZD.scala 39:21]
  wire  _T_472; // @[LZD.scala 39:30]
  wire  _T_473; // @[LZD.scala 39:27]
  wire  _T_474; // @[LZD.scala 39:25]
  wire [1:0] _T_475; // @[Cat.scala 29:58]
  wire  _T_476; // @[Shift.scala 12:21]
  wire  _T_477; // @[Shift.scala 12:21]
  wire  _T_478; // @[LZD.scala 49:16]
  wire  _T_479; // @[LZD.scala 49:27]
  wire  _T_480; // @[LZD.scala 49:25]
  wire  _T_481; // @[LZD.scala 49:47]
  wire  _T_482; // @[LZD.scala 49:59]
  wire  _T_483; // @[LZD.scala 49:35]
  wire [2:0] _T_485; // @[Cat.scala 29:58]
  wire  _T_486; // @[Shift.scala 12:21]
  wire  _T_487; // @[Shift.scala 12:21]
  wire  _T_488; // @[LZD.scala 49:16]
  wire  _T_489; // @[LZD.scala 49:27]
  wire  _T_490; // @[LZD.scala 49:25]
  wire [1:0] _T_491; // @[LZD.scala 49:47]
  wire [1:0] _T_492; // @[LZD.scala 49:59]
  wire [1:0] _T_493; // @[LZD.scala 49:35]
  wire [3:0] _T_495; // @[Cat.scala 29:58]
  wire [3:0] _T_496; // @[LZD.scala 44:32]
  wire [1:0] _T_497; // @[LZD.scala 43:32]
  wire  _T_498; // @[LZD.scala 39:14]
  wire  _T_499; // @[LZD.scala 39:21]
  wire  _T_500; // @[LZD.scala 39:30]
  wire  _T_501; // @[LZD.scala 39:27]
  wire  _T_502; // @[LZD.scala 39:25]
  wire [1:0] _T_503; // @[Cat.scala 29:58]
  wire [1:0] _T_504; // @[LZD.scala 44:32]
  wire  _T_505; // @[LZD.scala 39:14]
  wire  _T_506; // @[LZD.scala 39:21]
  wire  _T_507; // @[LZD.scala 39:30]
  wire  _T_508; // @[LZD.scala 39:27]
  wire  _T_509; // @[LZD.scala 39:25]
  wire [1:0] _T_510; // @[Cat.scala 29:58]
  wire  _T_511; // @[Shift.scala 12:21]
  wire  _T_512; // @[Shift.scala 12:21]
  wire  _T_513; // @[LZD.scala 49:16]
  wire  _T_514; // @[LZD.scala 49:27]
  wire  _T_515; // @[LZD.scala 49:25]
  wire  _T_516; // @[LZD.scala 49:47]
  wire  _T_517; // @[LZD.scala 49:59]
  wire  _T_518; // @[LZD.scala 49:35]
  wire [2:0] _T_520; // @[Cat.scala 29:58]
  wire  _T_521; // @[Shift.scala 12:21]
  wire [2:0] _T_523; // @[LZD.scala 55:32]
  wire [2:0] _T_524; // @[LZD.scala 55:20]
  wire [3:0] _T_525; // @[Cat.scala 29:58]
  wire  _T_526; // @[Shift.scala 12:21]
  wire [3:0] _T_528; // @[LZD.scala 55:32]
  wire [3:0] _T_529; // @[LZD.scala 55:20]
  wire [4:0] _T_530; // @[Cat.scala 29:58]
  wire [4:0] _T_531; // @[convert.scala 21:22]
  wire [26:0] _T_532; // @[convert.scala 22:36]
  wire  _T_533; // @[Shift.scala 16:24]
  wire  _T_535; // @[Shift.scala 12:21]
  wire [10:0] _T_536; // @[Shift.scala 64:52]
  wire [26:0] _T_538; // @[Cat.scala 29:58]
  wire [26:0] _T_539; // @[Shift.scala 64:27]
  wire [3:0] _T_540; // @[Shift.scala 66:70]
  wire  _T_541; // @[Shift.scala 12:21]
  wire [18:0] _T_542; // @[Shift.scala 64:52]
  wire [26:0] _T_544; // @[Cat.scala 29:58]
  wire [26:0] _T_545; // @[Shift.scala 64:27]
  wire [2:0] _T_546; // @[Shift.scala 66:70]
  wire  _T_547; // @[Shift.scala 12:21]
  wire [22:0] _T_548; // @[Shift.scala 64:52]
  wire [26:0] _T_550; // @[Cat.scala 29:58]
  wire [26:0] _T_551; // @[Shift.scala 64:27]
  wire [1:0] _T_552; // @[Shift.scala 66:70]
  wire  _T_553; // @[Shift.scala 12:21]
  wire [24:0] _T_554; // @[Shift.scala 64:52]
  wire [26:0] _T_556; // @[Cat.scala 29:58]
  wire [26:0] _T_557; // @[Shift.scala 64:27]
  wire  _T_558; // @[Shift.scala 66:70]
  wire [25:0] _T_560; // @[Shift.scala 64:52]
  wire [26:0] _T_561; // @[Cat.scala 29:58]
  wire [26:0] _T_562; // @[Shift.scala 64:27]
  wire [26:0] _T_563; // @[Shift.scala 16:10]
  wire [2:0] _T_564; // @[convert.scala 23:34]
  wire [23:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_566; // @[convert.scala 25:26]
  wire [4:0] _T_568; // @[convert.scala 25:42]
  wire [2:0] _T_571; // @[convert.scala 26:67]
  wire [2:0] _T_572; // @[convert.scala 26:51]
  wire [8:0] _T_573; // @[Cat.scala 29:58]
  wire [28:0] _T_575; // @[convert.scala 29:56]
  wire  _T_576; // @[convert.scala 29:60]
  wire  _T_577; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_580; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [8:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_589; // @[Bitwise.scala 71:12]
  wire  _T_590; // @[PositDivisionSqrt.scala 80:40]
  wire [27:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_592; // @[PositDivisionSqrt.scala 82:31]
  wire [27:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_595; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_596; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_597; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_598; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_599; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_600; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_601; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_602; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_603; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_604; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [9:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_607; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_608; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_609; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_610; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_611; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_612; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_613; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_614; // @[PositDivisionSqrt.scala 117:30]
  wire [4:0] _T_616; // @[PositDivisionSqrt.scala 119:26]
  wire [4:0] _T_617; // @[PositDivisionSqrt.scala 118:20]
  wire [4:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [4:0] _T_618; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_620; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_621; // @[PositDivisionSqrt.scala 123:27]
  wire [4:0] _T_623; // @[PositDivisionSqrt.scala 123:52]
  wire [4:0] _T_624; // @[PositDivisionSqrt.scala 123:20]
  wire [4:0] _T_625; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_627; // @[PositDivisionSqrt.scala 124:27]
  wire [4:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [4:0] _T_629; // @[PositDivisionSqrt.scala 123:64]
  wire [7:0] _T_630; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_632; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_633; // @[PositDivisionSqrt.scala 137:28]
  wire [31:0] _T_634; // @[PositDivisionSqrt.scala 146:22]
  wire [29:0] _T_635; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_636; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_637; // @[PositDivisionSqrt.scala 148:23]
  wire [27:0] _T_638; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_639; // @[PositDivisionSqrt.scala 149:23]
  wire [28:0] _T_640; // @[PositDivisionSqrt.scala 149:46]
  wire [27:0] _T_641; // @[PositDivisionSqrt.scala 149:56]
  wire [27:0] _T_642; // @[PositDivisionSqrt.scala 149:16]
  wire [27:0] _T_643; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_644; // @[PositDivisionSqrt.scala 150:17]
  wire [27:0] _T_645; // @[PositDivisionSqrt.scala 150:16]
  wire [27:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_647; // @[PositDivisionSqrt.scala 152:29]
  wire [27:0] _T_648; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_649; // @[PositDivisionSqrt.scala 153:29]
  wire [24:0] _T_650; // @[PositDivisionSqrt.scala 153:22]
  wire [27:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [27:0] _T_651; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_653; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_654; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_655; // @[PositDivisionSqrt.scala 154:57]
  wire [27:0] _T_658; // @[Cat.scala 29:58]
  wire [27:0] _T_659; // @[PositDivisionSqrt.scala 154:22]
  wire [27:0] _T_660; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_662; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_663; // @[PositDivisionSqrt.scala 156:79]
  wire [23:0] _T_665; // @[Bitwise.scala 71:12]
  wire [26:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [26:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [26:0] _T_666; // @[PositDivisionSqrt.scala 156:53]
  wire [27:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [27:0] _T_667; // @[PositDivisionSqrt.scala 155:51]
  wire [25:0] _T_668; // @[PositDivisionSqrt.scala 157:53]
  wire [27:0] _GEN_14; // @[PositDivisionSqrt.scala 156:85]
  wire [27:0] _T_669; // @[PositDivisionSqrt.scala 156:85]
  wire [27:0] _T_670; // @[PositDivisionSqrt.scala 155:22]
  wire [27:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_672; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_673; // @[PositDivisionSqrt.scala 162:40]
  wire [27:0] _T_676; // @[PositDivisionSqrt.scala 163:97]
  wire [27:0] _T_678; // @[PositDivisionSqrt.scala 164:97]
  wire [27:0] _T_679; // @[PositDivisionSqrt.scala 161:92]
  wire [28:0] _T_684; // @[PositDivisionSqrt.scala 168:98]
  wire [27:0] _T_685; // @[PositDivisionSqrt.scala 168:108]
  wire [27:0] _T_687; // @[PositDivisionSqrt.scala 168:112]
  wire [27:0] _T_691; // @[PositDivisionSqrt.scala 169:112]
  wire [27:0] _T_692; // @[PositDivisionSqrt.scala 166:26]
  wire [27:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_693; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_694; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_696; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_697; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_698; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_699; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_700; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_702; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_703; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_704; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_705; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_706; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_709; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_710; // @[PositDivisionSqrt.scala 187:28]
  wire [27:0] _T_713; // @[PositDivisionSqrt.scala 188:47]
  wire [27:0] _T_714; // @[PositDivisionSqrt.scala 188:18]
  wire [25:0] _T_716; // @[PositDivisionSqrt.scala 189:18]
  wire [27:0] _GEN_15; // @[PositDivisionSqrt.scala 188:72]
  wire [27:0] _T_717; // @[PositDivisionSqrt.scala 188:72]
  wire [27:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [27:0] _T_719; // @[PositDivisionSqrt.scala 190:47]
  wire [27:0] _T_720; // @[PositDivisionSqrt.scala 190:18]
  wire [27:0] _T_721; // @[PositDivisionSqrt.scala 189:72]
  wire [1:0] _T_723; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [27:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [27:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [23:0] _T_726; // @[PositDivisionSqrt.scala 200:97]
  wire [23:0] _T_727; // @[PositDivisionSqrt.scala 201:97]
  wire [23:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_728; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_729; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_730; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_732; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_733; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_734; // @[Cat.scala 29:58]
  wire [2:0] _T_735; // @[PositDivisionSqrt.scala 209:63]
  wire [9:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [9:0] _T_737; // @[PositDivisionSqrt.scala 209:31]
  wire [9:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [9:0] _T_739; // @[Mux.scala 87:16]
  wire [9:0] _T_740; // @[Mux.scala 87:16]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [8:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [8:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [2:0] _T_745; // @[convert.scala 46:61]
  wire [2:0] _T_746; // @[convert.scala 46:52]
  wire [2:0] _T_748; // @[convert.scala 46:42]
  wire [5:0] _T_749; // @[convert.scala 48:34]
  wire  _T_750; // @[convert.scala 49:36]
  wire [5:0] _T_752; // @[convert.scala 50:36]
  wire [5:0] _T_753; // @[convert.scala 50:36]
  wire [5:0] _T_754; // @[convert.scala 50:28]
  wire  _T_755; // @[convert.scala 51:31]
  wire  _T_756; // @[convert.scala 52:43]
  wire [31:0] _T_760; // @[Cat.scala 29:58]
  wire [5:0] _T_761; // @[Shift.scala 39:17]
  wire  _T_762; // @[Shift.scala 39:24]
  wire [4:0] _T_763; // @[Shift.scala 40:44]
  wire [15:0] _T_764; // @[Shift.scala 90:30]
  wire [15:0] _T_765; // @[Shift.scala 90:48]
  wire  _T_766; // @[Shift.scala 90:57]
  wire [15:0] _GEN_20; // @[Shift.scala 90:39]
  wire [15:0] _T_767; // @[Shift.scala 90:39]
  wire  _T_768; // @[Shift.scala 12:21]
  wire  _T_769; // @[Shift.scala 12:21]
  wire [15:0] _T_771; // @[Bitwise.scala 71:12]
  wire [31:0] _T_772; // @[Cat.scala 29:58]
  wire [31:0] _T_773; // @[Shift.scala 91:22]
  wire [3:0] _T_774; // @[Shift.scala 92:77]
  wire [23:0] _T_775; // @[Shift.scala 90:30]
  wire [7:0] _T_776; // @[Shift.scala 90:48]
  wire  _T_777; // @[Shift.scala 90:57]
  wire [23:0] _GEN_21; // @[Shift.scala 90:39]
  wire [23:0] _T_778; // @[Shift.scala 90:39]
  wire  _T_779; // @[Shift.scala 12:21]
  wire  _T_780; // @[Shift.scala 12:21]
  wire [7:0] _T_782; // @[Bitwise.scala 71:12]
  wire [31:0] _T_783; // @[Cat.scala 29:58]
  wire [31:0] _T_784; // @[Shift.scala 91:22]
  wire [2:0] _T_785; // @[Shift.scala 92:77]
  wire [27:0] _T_786; // @[Shift.scala 90:30]
  wire [3:0] _T_787; // @[Shift.scala 90:48]
  wire  _T_788; // @[Shift.scala 90:57]
  wire [27:0] _GEN_22; // @[Shift.scala 90:39]
  wire [27:0] _T_789; // @[Shift.scala 90:39]
  wire  _T_790; // @[Shift.scala 12:21]
  wire  _T_791; // @[Shift.scala 12:21]
  wire [3:0] _T_793; // @[Bitwise.scala 71:12]
  wire [31:0] _T_794; // @[Cat.scala 29:58]
  wire [31:0] _T_795; // @[Shift.scala 91:22]
  wire [1:0] _T_796; // @[Shift.scala 92:77]
  wire [29:0] _T_797; // @[Shift.scala 90:30]
  wire [1:0] _T_798; // @[Shift.scala 90:48]
  wire  _T_799; // @[Shift.scala 90:57]
  wire [29:0] _GEN_23; // @[Shift.scala 90:39]
  wire [29:0] _T_800; // @[Shift.scala 90:39]
  wire  _T_801; // @[Shift.scala 12:21]
  wire  _T_802; // @[Shift.scala 12:21]
  wire [1:0] _T_804; // @[Bitwise.scala 71:12]
  wire [31:0] _T_805; // @[Cat.scala 29:58]
  wire [31:0] _T_806; // @[Shift.scala 91:22]
  wire  _T_807; // @[Shift.scala 92:77]
  wire [30:0] _T_808; // @[Shift.scala 90:30]
  wire  _T_809; // @[Shift.scala 90:48]
  wire [30:0] _GEN_24; // @[Shift.scala 90:39]
  wire [30:0] _T_811; // @[Shift.scala 90:39]
  wire  _T_813; // @[Shift.scala 12:21]
  wire [31:0] _T_814; // @[Cat.scala 29:58]
  wire [31:0] _T_815; // @[Shift.scala 91:22]
  wire [31:0] _T_818; // @[Bitwise.scala 71:12]
  wire [31:0] _T_819; // @[Shift.scala 39:10]
  wire  _T_820; // @[convert.scala 55:31]
  wire  _T_821; // @[convert.scala 56:31]
  wire  _T_822; // @[convert.scala 57:31]
  wire  _T_823; // @[convert.scala 58:31]
  wire [28:0] _T_824; // @[convert.scala 59:69]
  wire  _T_825; // @[convert.scala 59:81]
  wire  _T_826; // @[convert.scala 59:50]
  wire  _T_828; // @[convert.scala 60:81]
  wire  _T_829; // @[convert.scala 61:44]
  wire  _T_830; // @[convert.scala 61:52]
  wire  _T_831; // @[convert.scala 61:36]
  wire  _T_832; // @[convert.scala 62:63]
  wire  _T_833; // @[convert.scala 62:103]
  wire  _T_834; // @[convert.scala 62:60]
  wire [28:0] _GEN_25; // @[convert.scala 63:56]
  wire [28:0] _T_837; // @[convert.scala 63:56]
  wire [29:0] _T_838; // @[Cat.scala 29:58]
  wire [29:0] _T_840; // @[Mux.scala 87:16]
  assign _T_1 = io_A[29]; // @[convert.scala 18:24]
  assign _T_2 = io_A[28]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[28:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[27:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[27:12]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[15:8]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[7:4]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9[3:2]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10 != 2'h0; // @[LZD.scala 39:14]
  assign _T_12 = _T_10[1]; // @[LZD.scala 39:21]
  assign _T_13 = _T_10[0]; // @[LZD.scala 39:30]
  assign _T_14 = ~ _T_13; // @[LZD.scala 39:27]
  assign _T_15 = _T_12 | _T_14; // @[LZD.scala 39:25]
  assign _T_16 = {_T_11,_T_15}; // @[Cat.scala 29:58]
  assign _T_17 = _T_9[1:0]; // @[LZD.scala 44:32]
  assign _T_18 = _T_17 != 2'h0; // @[LZD.scala 39:14]
  assign _T_19 = _T_17[1]; // @[LZD.scala 39:21]
  assign _T_20 = _T_17[0]; // @[LZD.scala 39:30]
  assign _T_21 = ~ _T_20; // @[LZD.scala 39:27]
  assign _T_22 = _T_19 | _T_21; // @[LZD.scala 39:25]
  assign _T_23 = {_T_18,_T_22}; // @[Cat.scala 29:58]
  assign _T_24 = _T_16[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23[1]; // @[Shift.scala 12:21]
  assign _T_26 = _T_24 | _T_25; // @[LZD.scala 49:16]
  assign _T_27 = ~ _T_25; // @[LZD.scala 49:27]
  assign _T_28 = _T_24 | _T_27; // @[LZD.scala 49:25]
  assign _T_29 = _T_16[0:0]; // @[LZD.scala 49:47]
  assign _T_30 = _T_23[0:0]; // @[LZD.scala 49:59]
  assign _T_31 = _T_24 ? _T_29 : _T_30; // @[LZD.scala 49:35]
  assign _T_33 = {_T_26,_T_28,_T_31}; // @[Cat.scala 29:58]
  assign _T_34 = _T_8[3:0]; // @[LZD.scala 44:32]
  assign _T_35 = _T_34[3:2]; // @[LZD.scala 43:32]
  assign _T_36 = _T_35 != 2'h0; // @[LZD.scala 39:14]
  assign _T_37 = _T_35[1]; // @[LZD.scala 39:21]
  assign _T_38 = _T_35[0]; // @[LZD.scala 39:30]
  assign _T_39 = ~ _T_38; // @[LZD.scala 39:27]
  assign _T_40 = _T_37 | _T_39; // @[LZD.scala 39:25]
  assign _T_41 = {_T_36,_T_40}; // @[Cat.scala 29:58]
  assign _T_42 = _T_34[1:0]; // @[LZD.scala 44:32]
  assign _T_43 = _T_42 != 2'h0; // @[LZD.scala 39:14]
  assign _T_44 = _T_42[1]; // @[LZD.scala 39:21]
  assign _T_45 = _T_42[0]; // @[LZD.scala 39:30]
  assign _T_46 = ~ _T_45; // @[LZD.scala 39:27]
  assign _T_47 = _T_44 | _T_46; // @[LZD.scala 39:25]
  assign _T_48 = {_T_43,_T_47}; // @[Cat.scala 29:58]
  assign _T_49 = _T_41[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48[1]; // @[Shift.scala 12:21]
  assign _T_51 = _T_49 | _T_50; // @[LZD.scala 49:16]
  assign _T_52 = ~ _T_50; // @[LZD.scala 49:27]
  assign _T_53 = _T_49 | _T_52; // @[LZD.scala 49:25]
  assign _T_54 = _T_41[0:0]; // @[LZD.scala 49:47]
  assign _T_55 = _T_48[0:0]; // @[LZD.scala 49:59]
  assign _T_56 = _T_49 ? _T_54 : _T_55; // @[LZD.scala 49:35]
  assign _T_58 = {_T_51,_T_53,_T_56}; // @[Cat.scala 29:58]
  assign _T_59 = _T_33[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58[2]; // @[Shift.scala 12:21]
  assign _T_61 = _T_59 | _T_60; // @[LZD.scala 49:16]
  assign _T_62 = ~ _T_60; // @[LZD.scala 49:27]
  assign _T_63 = _T_59 | _T_62; // @[LZD.scala 49:25]
  assign _T_64 = _T_33[1:0]; // @[LZD.scala 49:47]
  assign _T_65 = _T_58[1:0]; // @[LZD.scala 49:59]
  assign _T_66 = _T_59 ? _T_64 : _T_65; // @[LZD.scala 49:35]
  assign _T_68 = {_T_61,_T_63,_T_66}; // @[Cat.scala 29:58]
  assign _T_69 = _T_7[7:0]; // @[LZD.scala 44:32]
  assign _T_70 = _T_69[7:4]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70[3:2]; // @[LZD.scala 43:32]
  assign _T_72 = _T_71 != 2'h0; // @[LZD.scala 39:14]
  assign _T_73 = _T_71[1]; // @[LZD.scala 39:21]
  assign _T_74 = _T_71[0]; // @[LZD.scala 39:30]
  assign _T_75 = ~ _T_74; // @[LZD.scala 39:27]
  assign _T_76 = _T_73 | _T_75; // @[LZD.scala 39:25]
  assign _T_77 = {_T_72,_T_76}; // @[Cat.scala 29:58]
  assign _T_78 = _T_70[1:0]; // @[LZD.scala 44:32]
  assign _T_79 = _T_78 != 2'h0; // @[LZD.scala 39:14]
  assign _T_80 = _T_78[1]; // @[LZD.scala 39:21]
  assign _T_81 = _T_78[0]; // @[LZD.scala 39:30]
  assign _T_82 = ~ _T_81; // @[LZD.scala 39:27]
  assign _T_83 = _T_80 | _T_82; // @[LZD.scala 39:25]
  assign _T_84 = {_T_79,_T_83}; // @[Cat.scala 29:58]
  assign _T_85 = _T_77[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84[1]; // @[Shift.scala 12:21]
  assign _T_87 = _T_85 | _T_86; // @[LZD.scala 49:16]
  assign _T_88 = ~ _T_86; // @[LZD.scala 49:27]
  assign _T_89 = _T_85 | _T_88; // @[LZD.scala 49:25]
  assign _T_90 = _T_77[0:0]; // @[LZD.scala 49:47]
  assign _T_91 = _T_84[0:0]; // @[LZD.scala 49:59]
  assign _T_92 = _T_85 ? _T_90 : _T_91; // @[LZD.scala 49:35]
  assign _T_94 = {_T_87,_T_89,_T_92}; // @[Cat.scala 29:58]
  assign _T_95 = _T_69[3:0]; // @[LZD.scala 44:32]
  assign _T_96 = _T_95[3:2]; // @[LZD.scala 43:32]
  assign _T_97 = _T_96 != 2'h0; // @[LZD.scala 39:14]
  assign _T_98 = _T_96[1]; // @[LZD.scala 39:21]
  assign _T_99 = _T_96[0]; // @[LZD.scala 39:30]
  assign _T_100 = ~ _T_99; // @[LZD.scala 39:27]
  assign _T_101 = _T_98 | _T_100; // @[LZD.scala 39:25]
  assign _T_102 = {_T_97,_T_101}; // @[Cat.scala 29:58]
  assign _T_103 = _T_95[1:0]; // @[LZD.scala 44:32]
  assign _T_104 = _T_103 != 2'h0; // @[LZD.scala 39:14]
  assign _T_105 = _T_103[1]; // @[LZD.scala 39:21]
  assign _T_106 = _T_103[0]; // @[LZD.scala 39:30]
  assign _T_107 = ~ _T_106; // @[LZD.scala 39:27]
  assign _T_108 = _T_105 | _T_107; // @[LZD.scala 39:25]
  assign _T_109 = {_T_104,_T_108}; // @[Cat.scala 29:58]
  assign _T_110 = _T_102[1]; // @[Shift.scala 12:21]
  assign _T_111 = _T_109[1]; // @[Shift.scala 12:21]
  assign _T_112 = _T_110 | _T_111; // @[LZD.scala 49:16]
  assign _T_113 = ~ _T_111; // @[LZD.scala 49:27]
  assign _T_114 = _T_110 | _T_113; // @[LZD.scala 49:25]
  assign _T_115 = _T_102[0:0]; // @[LZD.scala 49:47]
  assign _T_116 = _T_109[0:0]; // @[LZD.scala 49:59]
  assign _T_117 = _T_110 ? _T_115 : _T_116; // @[LZD.scala 49:35]
  assign _T_119 = {_T_112,_T_114,_T_117}; // @[Cat.scala 29:58]
  assign _T_120 = _T_94[2]; // @[Shift.scala 12:21]
  assign _T_121 = _T_119[2]; // @[Shift.scala 12:21]
  assign _T_122 = _T_120 | _T_121; // @[LZD.scala 49:16]
  assign _T_123 = ~ _T_121; // @[LZD.scala 49:27]
  assign _T_124 = _T_120 | _T_123; // @[LZD.scala 49:25]
  assign _T_125 = _T_94[1:0]; // @[LZD.scala 49:47]
  assign _T_126 = _T_119[1:0]; // @[LZD.scala 49:59]
  assign _T_127 = _T_120 ? _T_125 : _T_126; // @[LZD.scala 49:35]
  assign _T_129 = {_T_122,_T_124,_T_127}; // @[Cat.scala 29:58]
  assign _T_130 = _T_68[3]; // @[Shift.scala 12:21]
  assign _T_131 = _T_129[3]; // @[Shift.scala 12:21]
  assign _T_132 = _T_130 | _T_131; // @[LZD.scala 49:16]
  assign _T_133 = ~ _T_131; // @[LZD.scala 49:27]
  assign _T_134 = _T_130 | _T_133; // @[LZD.scala 49:25]
  assign _T_135 = _T_68[2:0]; // @[LZD.scala 49:47]
  assign _T_136 = _T_129[2:0]; // @[LZD.scala 49:59]
  assign _T_137 = _T_130 ? _T_135 : _T_136; // @[LZD.scala 49:35]
  assign _T_139 = {_T_132,_T_134,_T_137}; // @[Cat.scala 29:58]
  assign _T_140 = _T_6[11:0]; // @[LZD.scala 44:32]
  assign _T_141 = _T_140[11:4]; // @[LZD.scala 43:32]
  assign _T_142 = _T_141[7:4]; // @[LZD.scala 43:32]
  assign _T_143 = _T_142[3:2]; // @[LZD.scala 43:32]
  assign _T_144 = _T_143 != 2'h0; // @[LZD.scala 39:14]
  assign _T_145 = _T_143[1]; // @[LZD.scala 39:21]
  assign _T_146 = _T_143[0]; // @[LZD.scala 39:30]
  assign _T_147 = ~ _T_146; // @[LZD.scala 39:27]
  assign _T_148 = _T_145 | _T_147; // @[LZD.scala 39:25]
  assign _T_149 = {_T_144,_T_148}; // @[Cat.scala 29:58]
  assign _T_150 = _T_142[1:0]; // @[LZD.scala 44:32]
  assign _T_151 = _T_150 != 2'h0; // @[LZD.scala 39:14]
  assign _T_152 = _T_150[1]; // @[LZD.scala 39:21]
  assign _T_153 = _T_150[0]; // @[LZD.scala 39:30]
  assign _T_154 = ~ _T_153; // @[LZD.scala 39:27]
  assign _T_155 = _T_152 | _T_154; // @[LZD.scala 39:25]
  assign _T_156 = {_T_151,_T_155}; // @[Cat.scala 29:58]
  assign _T_157 = _T_149[1]; // @[Shift.scala 12:21]
  assign _T_158 = _T_156[1]; // @[Shift.scala 12:21]
  assign _T_159 = _T_157 | _T_158; // @[LZD.scala 49:16]
  assign _T_160 = ~ _T_158; // @[LZD.scala 49:27]
  assign _T_161 = _T_157 | _T_160; // @[LZD.scala 49:25]
  assign _T_162 = _T_149[0:0]; // @[LZD.scala 49:47]
  assign _T_163 = _T_156[0:0]; // @[LZD.scala 49:59]
  assign _T_164 = _T_157 ? _T_162 : _T_163; // @[LZD.scala 49:35]
  assign _T_166 = {_T_159,_T_161,_T_164}; // @[Cat.scala 29:58]
  assign _T_167 = _T_141[3:0]; // @[LZD.scala 44:32]
  assign _T_168 = _T_167[3:2]; // @[LZD.scala 43:32]
  assign _T_169 = _T_168 != 2'h0; // @[LZD.scala 39:14]
  assign _T_170 = _T_168[1]; // @[LZD.scala 39:21]
  assign _T_171 = _T_168[0]; // @[LZD.scala 39:30]
  assign _T_172 = ~ _T_171; // @[LZD.scala 39:27]
  assign _T_173 = _T_170 | _T_172; // @[LZD.scala 39:25]
  assign _T_174 = {_T_169,_T_173}; // @[Cat.scala 29:58]
  assign _T_175 = _T_167[1:0]; // @[LZD.scala 44:32]
  assign _T_176 = _T_175 != 2'h0; // @[LZD.scala 39:14]
  assign _T_177 = _T_175[1]; // @[LZD.scala 39:21]
  assign _T_178 = _T_175[0]; // @[LZD.scala 39:30]
  assign _T_179 = ~ _T_178; // @[LZD.scala 39:27]
  assign _T_180 = _T_177 | _T_179; // @[LZD.scala 39:25]
  assign _T_181 = {_T_176,_T_180}; // @[Cat.scala 29:58]
  assign _T_182 = _T_174[1]; // @[Shift.scala 12:21]
  assign _T_183 = _T_181[1]; // @[Shift.scala 12:21]
  assign _T_184 = _T_182 | _T_183; // @[LZD.scala 49:16]
  assign _T_185 = ~ _T_183; // @[LZD.scala 49:27]
  assign _T_186 = _T_182 | _T_185; // @[LZD.scala 49:25]
  assign _T_187 = _T_174[0:0]; // @[LZD.scala 49:47]
  assign _T_188 = _T_181[0:0]; // @[LZD.scala 49:59]
  assign _T_189 = _T_182 ? _T_187 : _T_188; // @[LZD.scala 49:35]
  assign _T_191 = {_T_184,_T_186,_T_189}; // @[Cat.scala 29:58]
  assign _T_192 = _T_166[2]; // @[Shift.scala 12:21]
  assign _T_193 = _T_191[2]; // @[Shift.scala 12:21]
  assign _T_194 = _T_192 | _T_193; // @[LZD.scala 49:16]
  assign _T_195 = ~ _T_193; // @[LZD.scala 49:27]
  assign _T_196 = _T_192 | _T_195; // @[LZD.scala 49:25]
  assign _T_197 = _T_166[1:0]; // @[LZD.scala 49:47]
  assign _T_198 = _T_191[1:0]; // @[LZD.scala 49:59]
  assign _T_199 = _T_192 ? _T_197 : _T_198; // @[LZD.scala 49:35]
  assign _T_201 = {_T_194,_T_196,_T_199}; // @[Cat.scala 29:58]
  assign _T_202 = _T_140[3:0]; // @[LZD.scala 44:32]
  assign _T_203 = _T_202[3:2]; // @[LZD.scala 43:32]
  assign _T_204 = _T_203 != 2'h0; // @[LZD.scala 39:14]
  assign _T_205 = _T_203[1]; // @[LZD.scala 39:21]
  assign _T_206 = _T_203[0]; // @[LZD.scala 39:30]
  assign _T_207 = ~ _T_206; // @[LZD.scala 39:27]
  assign _T_208 = _T_205 | _T_207; // @[LZD.scala 39:25]
  assign _T_209 = {_T_204,_T_208}; // @[Cat.scala 29:58]
  assign _T_210 = _T_202[1:0]; // @[LZD.scala 44:32]
  assign _T_211 = _T_210 != 2'h0; // @[LZD.scala 39:14]
  assign _T_212 = _T_210[1]; // @[LZD.scala 39:21]
  assign _T_213 = _T_210[0]; // @[LZD.scala 39:30]
  assign _T_214 = ~ _T_213; // @[LZD.scala 39:27]
  assign _T_215 = _T_212 | _T_214; // @[LZD.scala 39:25]
  assign _T_216 = {_T_211,_T_215}; // @[Cat.scala 29:58]
  assign _T_217 = _T_209[1]; // @[Shift.scala 12:21]
  assign _T_218 = _T_216[1]; // @[Shift.scala 12:21]
  assign _T_219 = _T_217 | _T_218; // @[LZD.scala 49:16]
  assign _T_220 = ~ _T_218; // @[LZD.scala 49:27]
  assign _T_221 = _T_217 | _T_220; // @[LZD.scala 49:25]
  assign _T_222 = _T_209[0:0]; // @[LZD.scala 49:47]
  assign _T_223 = _T_216[0:0]; // @[LZD.scala 49:59]
  assign _T_224 = _T_217 ? _T_222 : _T_223; // @[LZD.scala 49:35]
  assign _T_226 = {_T_219,_T_221,_T_224}; // @[Cat.scala 29:58]
  assign _T_227 = _T_201[3]; // @[Shift.scala 12:21]
  assign _T_229 = _T_201[2:0]; // @[LZD.scala 55:32]
  assign _T_230 = _T_227 ? _T_229 : _T_226; // @[LZD.scala 55:20]
  assign _T_231 = {_T_227,_T_230}; // @[Cat.scala 29:58]
  assign _T_232 = _T_139[4]; // @[Shift.scala 12:21]
  assign _T_234 = _T_139[3:0]; // @[LZD.scala 55:32]
  assign _T_235 = _T_232 ? _T_234 : _T_231; // @[LZD.scala 55:20]
  assign _T_236 = {_T_232,_T_235}; // @[Cat.scala 29:58]
  assign _T_237 = ~ _T_236; // @[convert.scala 21:22]
  assign _T_238 = io_A[26:0]; // @[convert.scala 22:36]
  assign _T_239 = _T_237 < 5'h1b; // @[Shift.scala 16:24]
  assign _T_241 = _T_237[4]; // @[Shift.scala 12:21]
  assign _T_242 = _T_238[10:0]; // @[Shift.scala 64:52]
  assign _T_244 = {_T_242,16'h0}; // @[Cat.scala 29:58]
  assign _T_245 = _T_241 ? _T_244 : _T_238; // @[Shift.scala 64:27]
  assign _T_246 = _T_237[3:0]; // @[Shift.scala 66:70]
  assign _T_247 = _T_246[3]; // @[Shift.scala 12:21]
  assign _T_248 = _T_245[18:0]; // @[Shift.scala 64:52]
  assign _T_250 = {_T_248,8'h0}; // @[Cat.scala 29:58]
  assign _T_251 = _T_247 ? _T_250 : _T_245; // @[Shift.scala 64:27]
  assign _T_252 = _T_246[2:0]; // @[Shift.scala 66:70]
  assign _T_253 = _T_252[2]; // @[Shift.scala 12:21]
  assign _T_254 = _T_251[22:0]; // @[Shift.scala 64:52]
  assign _T_256 = {_T_254,4'h0}; // @[Cat.scala 29:58]
  assign _T_257 = _T_253 ? _T_256 : _T_251; // @[Shift.scala 64:27]
  assign _T_258 = _T_252[1:0]; // @[Shift.scala 66:70]
  assign _T_259 = _T_258[1]; // @[Shift.scala 12:21]
  assign _T_260 = _T_257[24:0]; // @[Shift.scala 64:52]
  assign _T_262 = {_T_260,2'h0}; // @[Cat.scala 29:58]
  assign _T_263 = _T_259 ? _T_262 : _T_257; // @[Shift.scala 64:27]
  assign _T_264 = _T_258[0:0]; // @[Shift.scala 66:70]
  assign _T_266 = _T_263[25:0]; // @[Shift.scala 64:52]
  assign _T_267 = {_T_266,1'h0}; // @[Cat.scala 29:58]
  assign _T_268 = _T_264 ? _T_267 : _T_263; // @[Shift.scala 64:27]
  assign _T_269 = _T_239 ? _T_268 : 27'h0; // @[Shift.scala 16:10]
  assign _T_270 = _T_269[26:24]; // @[convert.scala 23:34]
  assign decA_fraction = _T_269[23:0]; // @[convert.scala 24:34]
  assign _T_272 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_274 = _T_3 ? _T_237 : _T_236; // @[convert.scala 25:42]
  assign _T_277 = ~ _T_270; // @[convert.scala 26:67]
  assign _T_278 = _T_1 ? _T_277 : _T_270; // @[convert.scala 26:51]
  assign _T_279 = {_T_272,_T_274,_T_278}; // @[Cat.scala 29:58]
  assign _T_281 = io_A[28:0]; // @[convert.scala 29:56]
  assign _T_282 = _T_281 != 29'h0; // @[convert.scala 29:60]
  assign _T_283 = ~ _T_282; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_283; // @[convert.scala 29:39]
  assign _T_286 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_286 & _T_283; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_279); // @[convert.scala 32:24]
  assign _T_295 = io_B[29]; // @[convert.scala 18:24]
  assign _T_296 = io_B[28]; // @[convert.scala 18:40]
  assign _T_297 = _T_295 ^ _T_296; // @[convert.scala 18:36]
  assign _T_298 = io_B[28:1]; // @[convert.scala 19:24]
  assign _T_299 = io_B[27:0]; // @[convert.scala 19:43]
  assign _T_300 = _T_298 ^ _T_299; // @[convert.scala 19:39]
  assign _T_301 = _T_300[27:12]; // @[LZD.scala 43:32]
  assign _T_302 = _T_301[15:8]; // @[LZD.scala 43:32]
  assign _T_303 = _T_302[7:4]; // @[LZD.scala 43:32]
  assign _T_304 = _T_303[3:2]; // @[LZD.scala 43:32]
  assign _T_305 = _T_304 != 2'h0; // @[LZD.scala 39:14]
  assign _T_306 = _T_304[1]; // @[LZD.scala 39:21]
  assign _T_307 = _T_304[0]; // @[LZD.scala 39:30]
  assign _T_308 = ~ _T_307; // @[LZD.scala 39:27]
  assign _T_309 = _T_306 | _T_308; // @[LZD.scala 39:25]
  assign _T_310 = {_T_305,_T_309}; // @[Cat.scala 29:58]
  assign _T_311 = _T_303[1:0]; // @[LZD.scala 44:32]
  assign _T_312 = _T_311 != 2'h0; // @[LZD.scala 39:14]
  assign _T_313 = _T_311[1]; // @[LZD.scala 39:21]
  assign _T_314 = _T_311[0]; // @[LZD.scala 39:30]
  assign _T_315 = ~ _T_314; // @[LZD.scala 39:27]
  assign _T_316 = _T_313 | _T_315; // @[LZD.scala 39:25]
  assign _T_317 = {_T_312,_T_316}; // @[Cat.scala 29:58]
  assign _T_318 = _T_310[1]; // @[Shift.scala 12:21]
  assign _T_319 = _T_317[1]; // @[Shift.scala 12:21]
  assign _T_320 = _T_318 | _T_319; // @[LZD.scala 49:16]
  assign _T_321 = ~ _T_319; // @[LZD.scala 49:27]
  assign _T_322 = _T_318 | _T_321; // @[LZD.scala 49:25]
  assign _T_323 = _T_310[0:0]; // @[LZD.scala 49:47]
  assign _T_324 = _T_317[0:0]; // @[LZD.scala 49:59]
  assign _T_325 = _T_318 ? _T_323 : _T_324; // @[LZD.scala 49:35]
  assign _T_327 = {_T_320,_T_322,_T_325}; // @[Cat.scala 29:58]
  assign _T_328 = _T_302[3:0]; // @[LZD.scala 44:32]
  assign _T_329 = _T_328[3:2]; // @[LZD.scala 43:32]
  assign _T_330 = _T_329 != 2'h0; // @[LZD.scala 39:14]
  assign _T_331 = _T_329[1]; // @[LZD.scala 39:21]
  assign _T_332 = _T_329[0]; // @[LZD.scala 39:30]
  assign _T_333 = ~ _T_332; // @[LZD.scala 39:27]
  assign _T_334 = _T_331 | _T_333; // @[LZD.scala 39:25]
  assign _T_335 = {_T_330,_T_334}; // @[Cat.scala 29:58]
  assign _T_336 = _T_328[1:0]; // @[LZD.scala 44:32]
  assign _T_337 = _T_336 != 2'h0; // @[LZD.scala 39:14]
  assign _T_338 = _T_336[1]; // @[LZD.scala 39:21]
  assign _T_339 = _T_336[0]; // @[LZD.scala 39:30]
  assign _T_340 = ~ _T_339; // @[LZD.scala 39:27]
  assign _T_341 = _T_338 | _T_340; // @[LZD.scala 39:25]
  assign _T_342 = {_T_337,_T_341}; // @[Cat.scala 29:58]
  assign _T_343 = _T_335[1]; // @[Shift.scala 12:21]
  assign _T_344 = _T_342[1]; // @[Shift.scala 12:21]
  assign _T_345 = _T_343 | _T_344; // @[LZD.scala 49:16]
  assign _T_346 = ~ _T_344; // @[LZD.scala 49:27]
  assign _T_347 = _T_343 | _T_346; // @[LZD.scala 49:25]
  assign _T_348 = _T_335[0:0]; // @[LZD.scala 49:47]
  assign _T_349 = _T_342[0:0]; // @[LZD.scala 49:59]
  assign _T_350 = _T_343 ? _T_348 : _T_349; // @[LZD.scala 49:35]
  assign _T_352 = {_T_345,_T_347,_T_350}; // @[Cat.scala 29:58]
  assign _T_353 = _T_327[2]; // @[Shift.scala 12:21]
  assign _T_354 = _T_352[2]; // @[Shift.scala 12:21]
  assign _T_355 = _T_353 | _T_354; // @[LZD.scala 49:16]
  assign _T_356 = ~ _T_354; // @[LZD.scala 49:27]
  assign _T_357 = _T_353 | _T_356; // @[LZD.scala 49:25]
  assign _T_358 = _T_327[1:0]; // @[LZD.scala 49:47]
  assign _T_359 = _T_352[1:0]; // @[LZD.scala 49:59]
  assign _T_360 = _T_353 ? _T_358 : _T_359; // @[LZD.scala 49:35]
  assign _T_362 = {_T_355,_T_357,_T_360}; // @[Cat.scala 29:58]
  assign _T_363 = _T_301[7:0]; // @[LZD.scala 44:32]
  assign _T_364 = _T_363[7:4]; // @[LZD.scala 43:32]
  assign _T_365 = _T_364[3:2]; // @[LZD.scala 43:32]
  assign _T_366 = _T_365 != 2'h0; // @[LZD.scala 39:14]
  assign _T_367 = _T_365[1]; // @[LZD.scala 39:21]
  assign _T_368 = _T_365[0]; // @[LZD.scala 39:30]
  assign _T_369 = ~ _T_368; // @[LZD.scala 39:27]
  assign _T_370 = _T_367 | _T_369; // @[LZD.scala 39:25]
  assign _T_371 = {_T_366,_T_370}; // @[Cat.scala 29:58]
  assign _T_372 = _T_364[1:0]; // @[LZD.scala 44:32]
  assign _T_373 = _T_372 != 2'h0; // @[LZD.scala 39:14]
  assign _T_374 = _T_372[1]; // @[LZD.scala 39:21]
  assign _T_375 = _T_372[0]; // @[LZD.scala 39:30]
  assign _T_376 = ~ _T_375; // @[LZD.scala 39:27]
  assign _T_377 = _T_374 | _T_376; // @[LZD.scala 39:25]
  assign _T_378 = {_T_373,_T_377}; // @[Cat.scala 29:58]
  assign _T_379 = _T_371[1]; // @[Shift.scala 12:21]
  assign _T_380 = _T_378[1]; // @[Shift.scala 12:21]
  assign _T_381 = _T_379 | _T_380; // @[LZD.scala 49:16]
  assign _T_382 = ~ _T_380; // @[LZD.scala 49:27]
  assign _T_383 = _T_379 | _T_382; // @[LZD.scala 49:25]
  assign _T_384 = _T_371[0:0]; // @[LZD.scala 49:47]
  assign _T_385 = _T_378[0:0]; // @[LZD.scala 49:59]
  assign _T_386 = _T_379 ? _T_384 : _T_385; // @[LZD.scala 49:35]
  assign _T_388 = {_T_381,_T_383,_T_386}; // @[Cat.scala 29:58]
  assign _T_389 = _T_363[3:0]; // @[LZD.scala 44:32]
  assign _T_390 = _T_389[3:2]; // @[LZD.scala 43:32]
  assign _T_391 = _T_390 != 2'h0; // @[LZD.scala 39:14]
  assign _T_392 = _T_390[1]; // @[LZD.scala 39:21]
  assign _T_393 = _T_390[0]; // @[LZD.scala 39:30]
  assign _T_394 = ~ _T_393; // @[LZD.scala 39:27]
  assign _T_395 = _T_392 | _T_394; // @[LZD.scala 39:25]
  assign _T_396 = {_T_391,_T_395}; // @[Cat.scala 29:58]
  assign _T_397 = _T_389[1:0]; // @[LZD.scala 44:32]
  assign _T_398 = _T_397 != 2'h0; // @[LZD.scala 39:14]
  assign _T_399 = _T_397[1]; // @[LZD.scala 39:21]
  assign _T_400 = _T_397[0]; // @[LZD.scala 39:30]
  assign _T_401 = ~ _T_400; // @[LZD.scala 39:27]
  assign _T_402 = _T_399 | _T_401; // @[LZD.scala 39:25]
  assign _T_403 = {_T_398,_T_402}; // @[Cat.scala 29:58]
  assign _T_404 = _T_396[1]; // @[Shift.scala 12:21]
  assign _T_405 = _T_403[1]; // @[Shift.scala 12:21]
  assign _T_406 = _T_404 | _T_405; // @[LZD.scala 49:16]
  assign _T_407 = ~ _T_405; // @[LZD.scala 49:27]
  assign _T_408 = _T_404 | _T_407; // @[LZD.scala 49:25]
  assign _T_409 = _T_396[0:0]; // @[LZD.scala 49:47]
  assign _T_410 = _T_403[0:0]; // @[LZD.scala 49:59]
  assign _T_411 = _T_404 ? _T_409 : _T_410; // @[LZD.scala 49:35]
  assign _T_413 = {_T_406,_T_408,_T_411}; // @[Cat.scala 29:58]
  assign _T_414 = _T_388[2]; // @[Shift.scala 12:21]
  assign _T_415 = _T_413[2]; // @[Shift.scala 12:21]
  assign _T_416 = _T_414 | _T_415; // @[LZD.scala 49:16]
  assign _T_417 = ~ _T_415; // @[LZD.scala 49:27]
  assign _T_418 = _T_414 | _T_417; // @[LZD.scala 49:25]
  assign _T_419 = _T_388[1:0]; // @[LZD.scala 49:47]
  assign _T_420 = _T_413[1:0]; // @[LZD.scala 49:59]
  assign _T_421 = _T_414 ? _T_419 : _T_420; // @[LZD.scala 49:35]
  assign _T_423 = {_T_416,_T_418,_T_421}; // @[Cat.scala 29:58]
  assign _T_424 = _T_362[3]; // @[Shift.scala 12:21]
  assign _T_425 = _T_423[3]; // @[Shift.scala 12:21]
  assign _T_426 = _T_424 | _T_425; // @[LZD.scala 49:16]
  assign _T_427 = ~ _T_425; // @[LZD.scala 49:27]
  assign _T_428 = _T_424 | _T_427; // @[LZD.scala 49:25]
  assign _T_429 = _T_362[2:0]; // @[LZD.scala 49:47]
  assign _T_430 = _T_423[2:0]; // @[LZD.scala 49:59]
  assign _T_431 = _T_424 ? _T_429 : _T_430; // @[LZD.scala 49:35]
  assign _T_433 = {_T_426,_T_428,_T_431}; // @[Cat.scala 29:58]
  assign _T_434 = _T_300[11:0]; // @[LZD.scala 44:32]
  assign _T_435 = _T_434[11:4]; // @[LZD.scala 43:32]
  assign _T_436 = _T_435[7:4]; // @[LZD.scala 43:32]
  assign _T_437 = _T_436[3:2]; // @[LZD.scala 43:32]
  assign _T_438 = _T_437 != 2'h0; // @[LZD.scala 39:14]
  assign _T_439 = _T_437[1]; // @[LZD.scala 39:21]
  assign _T_440 = _T_437[0]; // @[LZD.scala 39:30]
  assign _T_441 = ~ _T_440; // @[LZD.scala 39:27]
  assign _T_442 = _T_439 | _T_441; // @[LZD.scala 39:25]
  assign _T_443 = {_T_438,_T_442}; // @[Cat.scala 29:58]
  assign _T_444 = _T_436[1:0]; // @[LZD.scala 44:32]
  assign _T_445 = _T_444 != 2'h0; // @[LZD.scala 39:14]
  assign _T_446 = _T_444[1]; // @[LZD.scala 39:21]
  assign _T_447 = _T_444[0]; // @[LZD.scala 39:30]
  assign _T_448 = ~ _T_447; // @[LZD.scala 39:27]
  assign _T_449 = _T_446 | _T_448; // @[LZD.scala 39:25]
  assign _T_450 = {_T_445,_T_449}; // @[Cat.scala 29:58]
  assign _T_451 = _T_443[1]; // @[Shift.scala 12:21]
  assign _T_452 = _T_450[1]; // @[Shift.scala 12:21]
  assign _T_453 = _T_451 | _T_452; // @[LZD.scala 49:16]
  assign _T_454 = ~ _T_452; // @[LZD.scala 49:27]
  assign _T_455 = _T_451 | _T_454; // @[LZD.scala 49:25]
  assign _T_456 = _T_443[0:0]; // @[LZD.scala 49:47]
  assign _T_457 = _T_450[0:0]; // @[LZD.scala 49:59]
  assign _T_458 = _T_451 ? _T_456 : _T_457; // @[LZD.scala 49:35]
  assign _T_460 = {_T_453,_T_455,_T_458}; // @[Cat.scala 29:58]
  assign _T_461 = _T_435[3:0]; // @[LZD.scala 44:32]
  assign _T_462 = _T_461[3:2]; // @[LZD.scala 43:32]
  assign _T_463 = _T_462 != 2'h0; // @[LZD.scala 39:14]
  assign _T_464 = _T_462[1]; // @[LZD.scala 39:21]
  assign _T_465 = _T_462[0]; // @[LZD.scala 39:30]
  assign _T_466 = ~ _T_465; // @[LZD.scala 39:27]
  assign _T_467 = _T_464 | _T_466; // @[LZD.scala 39:25]
  assign _T_468 = {_T_463,_T_467}; // @[Cat.scala 29:58]
  assign _T_469 = _T_461[1:0]; // @[LZD.scala 44:32]
  assign _T_470 = _T_469 != 2'h0; // @[LZD.scala 39:14]
  assign _T_471 = _T_469[1]; // @[LZD.scala 39:21]
  assign _T_472 = _T_469[0]; // @[LZD.scala 39:30]
  assign _T_473 = ~ _T_472; // @[LZD.scala 39:27]
  assign _T_474 = _T_471 | _T_473; // @[LZD.scala 39:25]
  assign _T_475 = {_T_470,_T_474}; // @[Cat.scala 29:58]
  assign _T_476 = _T_468[1]; // @[Shift.scala 12:21]
  assign _T_477 = _T_475[1]; // @[Shift.scala 12:21]
  assign _T_478 = _T_476 | _T_477; // @[LZD.scala 49:16]
  assign _T_479 = ~ _T_477; // @[LZD.scala 49:27]
  assign _T_480 = _T_476 | _T_479; // @[LZD.scala 49:25]
  assign _T_481 = _T_468[0:0]; // @[LZD.scala 49:47]
  assign _T_482 = _T_475[0:0]; // @[LZD.scala 49:59]
  assign _T_483 = _T_476 ? _T_481 : _T_482; // @[LZD.scala 49:35]
  assign _T_485 = {_T_478,_T_480,_T_483}; // @[Cat.scala 29:58]
  assign _T_486 = _T_460[2]; // @[Shift.scala 12:21]
  assign _T_487 = _T_485[2]; // @[Shift.scala 12:21]
  assign _T_488 = _T_486 | _T_487; // @[LZD.scala 49:16]
  assign _T_489 = ~ _T_487; // @[LZD.scala 49:27]
  assign _T_490 = _T_486 | _T_489; // @[LZD.scala 49:25]
  assign _T_491 = _T_460[1:0]; // @[LZD.scala 49:47]
  assign _T_492 = _T_485[1:0]; // @[LZD.scala 49:59]
  assign _T_493 = _T_486 ? _T_491 : _T_492; // @[LZD.scala 49:35]
  assign _T_495 = {_T_488,_T_490,_T_493}; // @[Cat.scala 29:58]
  assign _T_496 = _T_434[3:0]; // @[LZD.scala 44:32]
  assign _T_497 = _T_496[3:2]; // @[LZD.scala 43:32]
  assign _T_498 = _T_497 != 2'h0; // @[LZD.scala 39:14]
  assign _T_499 = _T_497[1]; // @[LZD.scala 39:21]
  assign _T_500 = _T_497[0]; // @[LZD.scala 39:30]
  assign _T_501 = ~ _T_500; // @[LZD.scala 39:27]
  assign _T_502 = _T_499 | _T_501; // @[LZD.scala 39:25]
  assign _T_503 = {_T_498,_T_502}; // @[Cat.scala 29:58]
  assign _T_504 = _T_496[1:0]; // @[LZD.scala 44:32]
  assign _T_505 = _T_504 != 2'h0; // @[LZD.scala 39:14]
  assign _T_506 = _T_504[1]; // @[LZD.scala 39:21]
  assign _T_507 = _T_504[0]; // @[LZD.scala 39:30]
  assign _T_508 = ~ _T_507; // @[LZD.scala 39:27]
  assign _T_509 = _T_506 | _T_508; // @[LZD.scala 39:25]
  assign _T_510 = {_T_505,_T_509}; // @[Cat.scala 29:58]
  assign _T_511 = _T_503[1]; // @[Shift.scala 12:21]
  assign _T_512 = _T_510[1]; // @[Shift.scala 12:21]
  assign _T_513 = _T_511 | _T_512; // @[LZD.scala 49:16]
  assign _T_514 = ~ _T_512; // @[LZD.scala 49:27]
  assign _T_515 = _T_511 | _T_514; // @[LZD.scala 49:25]
  assign _T_516 = _T_503[0:0]; // @[LZD.scala 49:47]
  assign _T_517 = _T_510[0:0]; // @[LZD.scala 49:59]
  assign _T_518 = _T_511 ? _T_516 : _T_517; // @[LZD.scala 49:35]
  assign _T_520 = {_T_513,_T_515,_T_518}; // @[Cat.scala 29:58]
  assign _T_521 = _T_495[3]; // @[Shift.scala 12:21]
  assign _T_523 = _T_495[2:0]; // @[LZD.scala 55:32]
  assign _T_524 = _T_521 ? _T_523 : _T_520; // @[LZD.scala 55:20]
  assign _T_525 = {_T_521,_T_524}; // @[Cat.scala 29:58]
  assign _T_526 = _T_433[4]; // @[Shift.scala 12:21]
  assign _T_528 = _T_433[3:0]; // @[LZD.scala 55:32]
  assign _T_529 = _T_526 ? _T_528 : _T_525; // @[LZD.scala 55:20]
  assign _T_530 = {_T_526,_T_529}; // @[Cat.scala 29:58]
  assign _T_531 = ~ _T_530; // @[convert.scala 21:22]
  assign _T_532 = io_B[26:0]; // @[convert.scala 22:36]
  assign _T_533 = _T_531 < 5'h1b; // @[Shift.scala 16:24]
  assign _T_535 = _T_531[4]; // @[Shift.scala 12:21]
  assign _T_536 = _T_532[10:0]; // @[Shift.scala 64:52]
  assign _T_538 = {_T_536,16'h0}; // @[Cat.scala 29:58]
  assign _T_539 = _T_535 ? _T_538 : _T_532; // @[Shift.scala 64:27]
  assign _T_540 = _T_531[3:0]; // @[Shift.scala 66:70]
  assign _T_541 = _T_540[3]; // @[Shift.scala 12:21]
  assign _T_542 = _T_539[18:0]; // @[Shift.scala 64:52]
  assign _T_544 = {_T_542,8'h0}; // @[Cat.scala 29:58]
  assign _T_545 = _T_541 ? _T_544 : _T_539; // @[Shift.scala 64:27]
  assign _T_546 = _T_540[2:0]; // @[Shift.scala 66:70]
  assign _T_547 = _T_546[2]; // @[Shift.scala 12:21]
  assign _T_548 = _T_545[22:0]; // @[Shift.scala 64:52]
  assign _T_550 = {_T_548,4'h0}; // @[Cat.scala 29:58]
  assign _T_551 = _T_547 ? _T_550 : _T_545; // @[Shift.scala 64:27]
  assign _T_552 = _T_546[1:0]; // @[Shift.scala 66:70]
  assign _T_553 = _T_552[1]; // @[Shift.scala 12:21]
  assign _T_554 = _T_551[24:0]; // @[Shift.scala 64:52]
  assign _T_556 = {_T_554,2'h0}; // @[Cat.scala 29:58]
  assign _T_557 = _T_553 ? _T_556 : _T_551; // @[Shift.scala 64:27]
  assign _T_558 = _T_552[0:0]; // @[Shift.scala 66:70]
  assign _T_560 = _T_557[25:0]; // @[Shift.scala 64:52]
  assign _T_561 = {_T_560,1'h0}; // @[Cat.scala 29:58]
  assign _T_562 = _T_558 ? _T_561 : _T_557; // @[Shift.scala 64:27]
  assign _T_563 = _T_533 ? _T_562 : 27'h0; // @[Shift.scala 16:10]
  assign _T_564 = _T_563[26:24]; // @[convert.scala 23:34]
  assign decB_fraction = _T_563[23:0]; // @[convert.scala 24:34]
  assign _T_566 = _T_297 == 1'h0; // @[convert.scala 25:26]
  assign _T_568 = _T_297 ? _T_531 : _T_530; // @[convert.scala 25:42]
  assign _T_571 = ~ _T_564; // @[convert.scala 26:67]
  assign _T_572 = _T_295 ? _T_571 : _T_564; // @[convert.scala 26:51]
  assign _T_573 = {_T_566,_T_568,_T_572}; // @[Cat.scala 29:58]
  assign _T_575 = io_B[28:0]; // @[convert.scala 29:56]
  assign _T_576 = _T_575 != 29'h0; // @[convert.scala 29:60]
  assign _T_577 = ~ _T_576; // @[convert.scala 29:41]
  assign decB_isNaR = _T_295 & _T_577; // @[convert.scala 29:39]
  assign _T_580 = _T_295 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_580 & _T_577; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_573); // @[convert.scala 32:24]
  assign _T_589 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_590 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_589,_T_590,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_592 = ~ _T_295; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_295,_T_592,decB_fraction,2'h0}; // @[Cat.scala 29:58]
  assign _T_595 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_595 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_596 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_597 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_598 = _T_597 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_599 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_600 = decA_isZero & _T_599; // @[PositDivisionSqrt.scala 94:43]
  assign _T_601 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_602 = _T_600 & _T_601; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_603 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_604 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_603 & _T_604; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_603 & _T_286; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_607 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_607; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 5'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 5'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_608 = sigX_Z[27]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_609 = sigX_Z[25]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_608 ^ _T_609; // @[PositDivisionSqrt.scala 113:50]
  assign _T_610 = cycleNum == 5'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_610 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_611 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_612 = _T_611 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_613 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_614 = entering & _T_613; // @[PositDivisionSqrt.scala 117:30]
  assign _T_616 = io_sqrtOp ? 5'h1a : 5'h1c; // @[PositDivisionSqrt.scala 119:26]
  assign _T_617 = entering_normalCase ? _T_616 : 5'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{4'd0}, _T_614}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_618 = _GEN_9 | _T_617; // @[PositDivisionSqrt.scala 117:64]
  assign _T_620 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_621 = _T_611 & _T_620; // @[PositDivisionSqrt.scala 123:27]
  assign _T_623 = cycleNum - 5'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_624 = _T_621 ? _T_623 : 5'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_625 = _T_618 | _T_624; // @[PositDivisionSqrt.scala 122:64]
  assign _T_627 = _T_611 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{4'd0}, _T_627}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_629 = _T_625 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_630 = decA_scale[8:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_632 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_633 = entering_normalCase & _T_632; // @[PositDivisionSqrt.scala 137:28]
  assign _T_634 = 32'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_635 = _T_634[31:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_636 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_637 = ready & _T_636; // @[PositDivisionSqrt.scala 148:23]
  assign _T_638 = _T_637 ? sigA_S : 28'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_639 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_640 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_641 = _T_640[27:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_642 = _T_639 ? _T_641 : 28'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_643 = _T_638 | _T_642; // @[PositDivisionSqrt.scala 148:66]
  assign _T_644 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_645 = _T_644 ? rem_Z : 28'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_643 | _T_645; // @[PositDivisionSqrt.scala 149:66]
  assign _T_647 = ready & _T_632; // @[PositDivisionSqrt.scala 152:29]
  assign _T_648 = _T_647 ? sigB_S : 28'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_649 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_650 = _T_649 ? 25'h1000000 : 25'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_650}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_651 = _T_648 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_653 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_654 = _T_644 & _T_653; // @[PositDivisionSqrt.scala 154:30]
  assign _T_655 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_658 = {signB_Z,_T_655,fractB_Z,2'h0}; // @[Cat.scala 29:58]
  assign _T_659 = _T_654 ? _T_658 : 28'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_660 = _T_651 | _T_659; // @[PositDivisionSqrt.scala 153:93]
  assign _T_662 = _T_644 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_663 = rem[27:27]; // @[PositDivisionSqrt.scala 156:79]
  assign _T_665 = _T_663 ? 24'hffffff : 24'h0; // @[Bitwise.scala 71:12]
  assign bitMask = _T_635[26:0]; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_12 = {{3'd0}, _T_665}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_666 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_666}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_667 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_668 = bitMask[26:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_668}; // @[PositDivisionSqrt.scala 156:85]
  assign _T_669 = _T_667 | _GEN_14; // @[PositDivisionSqrt.scala 156:85]
  assign _T_670 = _T_662 ? _T_669 : 28'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_660 | _T_670; // @[PositDivisionSqrt.scala 154:93]
  assign _T_672 = trialTerm[27:27]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_673 = _T_663 ^ _T_672; // @[PositDivisionSqrt.scala 162:40]
  assign _T_676 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_678 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_679 = _T_673 ? _T_676 : _T_678; // @[PositDivisionSqrt.scala 161:92]
  assign _T_684 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_685 = _T_684[27:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_687 = _T_685 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_691 = _T_685 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_692 = _T_673 ? _T_687 : _T_691; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_679 : _T_692; // @[PositDivisionSqrt.scala 159:27]
  assign _T_693 = trialRem != 28'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_693 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_694 = rem != 28'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_694 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_696 = trialRem[27:27]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_697 = _T_672 ^ _T_696; // @[PositDivisionSqrt.scala 176:49]
  assign _T_698 = ~ _T_697; // @[PositDivisionSqrt.scala 176:29]
  assign _T_699 = sigX_Z[27:27]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_700 = ~ _T_699; // @[PositDivisionSqrt.scala 178:49]
  assign _T_702 = remIsZero ? _T_699 : _T_698; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_700 : _T_702; // @[Mux.scala 87:16]
  assign _T_703 = cycleNum > 5'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_704 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_705 = _T_703 & _T_704; // @[PositDivisionSqrt.scala 183:48]
  assign _T_706 = entering_normalCase | _T_705; // @[PositDivisionSqrt.scala 183:28]
  assign _T_709 = _T_644 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_710 = entering_normalCase | _T_709; // @[PositDivisionSqrt.scala 187:28]
  assign _T_713 = {newBit, 27'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_714 = _T_647 ? _T_713 : 28'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_716 = _T_649 ? 26'h2000000 : 26'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_716}; // @[PositDivisionSqrt.scala 188:72]
  assign _T_717 = _T_714 | _GEN_15; // @[PositDivisionSqrt.scala 188:72]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_719 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_720 = _T_644 ? _T_719 : 28'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_721 = _T_717 | _T_720; // @[PositDivisionSqrt.scala 189:72]
  assign _T_723 = {_T_699, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_723 : {{1'd0}, _T_699}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{26'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_726 = realSigX[24:1]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_727 = realSigX[23:0]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_726 : _T_727; // @[PositDivisionSqrt.scala 198:21]
  assign _T_728 = realSigX[27]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_729 = realSigX[25]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_730 = _T_728 ^ _T_729; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_730; // @[PositDivisionSqrt.scala 205:23]
  assign _T_732 = realSigX[24]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_728 ^ _T_732; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_733 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_733; // @[PositDivisionSqrt.scala 208:36]
  assign _T_734 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_735 = {1'b0,$signed(_T_734)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{7{_T_735[2]}},_T_735}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_737 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_737); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-10'she0); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(10'she0); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[27:27]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_739 = underflow ? $signed(-10'she0) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_740 = overflow ? $signed(10'she0) : $signed(_T_739); // @[Mux.scala 87:16]
  assign outValid = cycleNum == 5'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_740[8:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_745 = decQ_scale[2:0]; // @[convert.scala 46:61]
  assign _T_746 = ~ _T_745; // @[convert.scala 46:52]
  assign _T_748 = decQ_sign ? _T_746 : _T_745; // @[convert.scala 46:42]
  assign _T_749 = decQ_scale[8:3]; // @[convert.scala 48:34]
  assign _T_750 = _T_749[5:5]; // @[convert.scala 49:36]
  assign _T_752 = ~ _T_749; // @[convert.scala 50:36]
  assign _T_753 = $signed(_T_752); // @[convert.scala 50:36]
  assign _T_754 = _T_750 ? $signed(_T_753) : $signed(_T_749); // @[convert.scala 50:28]
  assign _T_755 = _T_750 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_756 = ~ _T_755; // @[convert.scala 52:43]
  assign _T_760 = {_T_756,_T_755,_T_748,realFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_761 = $unsigned(_T_754); // @[Shift.scala 39:17]
  assign _T_762 = _T_761 < 6'h20; // @[Shift.scala 39:24]
  assign _T_763 = _T_754[4:0]; // @[Shift.scala 40:44]
  assign _T_764 = _T_760[31:16]; // @[Shift.scala 90:30]
  assign _T_765 = _T_760[15:0]; // @[Shift.scala 90:48]
  assign _T_766 = _T_765 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{15'd0}, _T_766}; // @[Shift.scala 90:39]
  assign _T_767 = _T_764 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_768 = _T_763[4]; // @[Shift.scala 12:21]
  assign _T_769 = _T_760[31]; // @[Shift.scala 12:21]
  assign _T_771 = _T_769 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_772 = {_T_771,_T_767}; // @[Cat.scala 29:58]
  assign _T_773 = _T_768 ? _T_772 : _T_760; // @[Shift.scala 91:22]
  assign _T_774 = _T_763[3:0]; // @[Shift.scala 92:77]
  assign _T_775 = _T_773[31:8]; // @[Shift.scala 90:30]
  assign _T_776 = _T_773[7:0]; // @[Shift.scala 90:48]
  assign _T_777 = _T_776 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{23'd0}, _T_777}; // @[Shift.scala 90:39]
  assign _T_778 = _T_775 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_779 = _T_774[3]; // @[Shift.scala 12:21]
  assign _T_780 = _T_773[31]; // @[Shift.scala 12:21]
  assign _T_782 = _T_780 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_783 = {_T_782,_T_778}; // @[Cat.scala 29:58]
  assign _T_784 = _T_779 ? _T_783 : _T_773; // @[Shift.scala 91:22]
  assign _T_785 = _T_774[2:0]; // @[Shift.scala 92:77]
  assign _T_786 = _T_784[31:4]; // @[Shift.scala 90:30]
  assign _T_787 = _T_784[3:0]; // @[Shift.scala 90:48]
  assign _T_788 = _T_787 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{27'd0}, _T_788}; // @[Shift.scala 90:39]
  assign _T_789 = _T_786 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_790 = _T_785[2]; // @[Shift.scala 12:21]
  assign _T_791 = _T_784[31]; // @[Shift.scala 12:21]
  assign _T_793 = _T_791 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_794 = {_T_793,_T_789}; // @[Cat.scala 29:58]
  assign _T_795 = _T_790 ? _T_794 : _T_784; // @[Shift.scala 91:22]
  assign _T_796 = _T_785[1:0]; // @[Shift.scala 92:77]
  assign _T_797 = _T_795[31:2]; // @[Shift.scala 90:30]
  assign _T_798 = _T_795[1:0]; // @[Shift.scala 90:48]
  assign _T_799 = _T_798 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{29'd0}, _T_799}; // @[Shift.scala 90:39]
  assign _T_800 = _T_797 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_801 = _T_796[1]; // @[Shift.scala 12:21]
  assign _T_802 = _T_795[31]; // @[Shift.scala 12:21]
  assign _T_804 = _T_802 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_805 = {_T_804,_T_800}; // @[Cat.scala 29:58]
  assign _T_806 = _T_801 ? _T_805 : _T_795; // @[Shift.scala 91:22]
  assign _T_807 = _T_796[0:0]; // @[Shift.scala 92:77]
  assign _T_808 = _T_806[31:1]; // @[Shift.scala 90:30]
  assign _T_809 = _T_806[0:0]; // @[Shift.scala 90:48]
  assign _GEN_24 = {{30'd0}, _T_809}; // @[Shift.scala 90:39]
  assign _T_811 = _T_808 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_813 = _T_806[31]; // @[Shift.scala 12:21]
  assign _T_814 = {_T_813,_T_811}; // @[Cat.scala 29:58]
  assign _T_815 = _T_807 ? _T_814 : _T_806; // @[Shift.scala 91:22]
  assign _T_818 = _T_769 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 71:12]
  assign _T_819 = _T_762 ? _T_815 : _T_818; // @[Shift.scala 39:10]
  assign _T_820 = _T_819[3]; // @[convert.scala 55:31]
  assign _T_821 = _T_819[2]; // @[convert.scala 56:31]
  assign _T_822 = _T_819[1]; // @[convert.scala 57:31]
  assign _T_823 = _T_819[0]; // @[convert.scala 58:31]
  assign _T_824 = _T_819[31:3]; // @[convert.scala 59:69]
  assign _T_825 = _T_824 != 29'h0; // @[convert.scala 59:81]
  assign _T_826 = ~ _T_825; // @[convert.scala 59:50]
  assign _T_828 = _T_824 == 29'h1fffffff; // @[convert.scala 60:81]
  assign _T_829 = _T_820 | _T_822; // @[convert.scala 61:44]
  assign _T_830 = _T_829 | _T_823; // @[convert.scala 61:52]
  assign _T_831 = _T_821 & _T_830; // @[convert.scala 61:36]
  assign _T_832 = ~ _T_828; // @[convert.scala 62:63]
  assign _T_833 = _T_832 & _T_831; // @[convert.scala 62:103]
  assign _T_834 = _T_826 | _T_833; // @[convert.scala 62:60]
  assign _GEN_25 = {{28'd0}, _T_834}; // @[convert.scala 63:56]
  assign _T_837 = _T_824 + _GEN_25; // @[convert.scala 63:56]
  assign _T_838 = {decQ_sign,_T_837}; // @[Cat.scala 29:58]
  assign _T_840 = isZero_Z ? 30'h0 : _T_838; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 5'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_653; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 30'h20000000 : _T_840; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[23:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[27:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[27:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 5'h0;
    end else begin
      if (_T_612) begin
        cycleNum <= _T_629;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_596;
      end else begin
        isNaR_Z <= _T_598;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_602;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_630[7]}},_T_630};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_633) begin
      signB_Z <= _T_295;
    end
    if (_T_633) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_706) begin
      if (ready) begin
        if (_T_673) begin
          rem_Z <= _T_676;
        end else begin
          rem_Z <= _T_678;
        end
      end else begin
        if (_T_673) begin
          rem_Z <= _T_687;
        end else begin
          rem_Z <= _T_691;
        end
      end
    end
    if (_T_710) begin
      sigX_Z <= _T_721;
    end
  end
endmodule
