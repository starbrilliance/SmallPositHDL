module PositAdder15_1(
  input         clock,
  input         reset,
  input  [14:0] io_A,
  input  [14:0] io_B,
  output [14:0] io_S
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [12:0] _T_4; // @[convert.scala 19:24]
  wire [12:0] _T_5; // @[convert.scala 19:43]
  wire [12:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [4:0] _T_68; // @[LZD.scala 44:32]
  wire [3:0] _T_69; // @[LZD.scala 43:32]
  wire [1:0] _T_70; // @[LZD.scala 43:32]
  wire  _T_71; // @[LZD.scala 39:14]
  wire  _T_72; // @[LZD.scala 39:21]
  wire  _T_73; // @[LZD.scala 39:30]
  wire  _T_74; // @[LZD.scala 39:27]
  wire  _T_75; // @[LZD.scala 39:25]
  wire [1:0] _T_76; // @[Cat.scala 29:58]
  wire [1:0] _T_77; // @[LZD.scala 44:32]
  wire  _T_78; // @[LZD.scala 39:14]
  wire  _T_79; // @[LZD.scala 39:21]
  wire  _T_80; // @[LZD.scala 39:30]
  wire  _T_81; // @[LZD.scala 39:27]
  wire  _T_82; // @[LZD.scala 39:25]
  wire [1:0] _T_83; // @[Cat.scala 29:58]
  wire  _T_84; // @[Shift.scala 12:21]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[LZD.scala 49:16]
  wire  _T_87; // @[LZD.scala 49:27]
  wire  _T_88; // @[LZD.scala 49:25]
  wire  _T_89; // @[LZD.scala 49:47]
  wire  _T_90; // @[LZD.scala 49:59]
  wire  _T_91; // @[LZD.scala 49:35]
  wire [2:0] _T_93; // @[Cat.scala 29:58]
  wire  _T_94; // @[LZD.scala 44:32]
  wire  _T_96; // @[Shift.scala 12:21]
  wire [1:0] _T_98; // @[Cat.scala 29:58]
  wire [1:0] _T_99; // @[LZD.scala 55:32]
  wire [1:0] _T_100; // @[LZD.scala 55:20]
  wire [2:0] _T_101; // @[Cat.scala 29:58]
  wire  _T_102; // @[Shift.scala 12:21]
  wire [2:0] _T_104; // @[LZD.scala 55:32]
  wire [2:0] _T_105; // @[LZD.scala 55:20]
  wire [3:0] _T_106; // @[Cat.scala 29:58]
  wire [3:0] _T_107; // @[convert.scala 21:22]
  wire [11:0] _T_108; // @[convert.scala 22:36]
  wire  _T_109; // @[Shift.scala 16:24]
  wire  _T_111; // @[Shift.scala 12:21]
  wire [3:0] _T_112; // @[Shift.scala 64:52]
  wire [11:0] _T_114; // @[Cat.scala 29:58]
  wire [11:0] _T_115; // @[Shift.scala 64:27]
  wire [2:0] _T_116; // @[Shift.scala 66:70]
  wire  _T_117; // @[Shift.scala 12:21]
  wire [7:0] _T_118; // @[Shift.scala 64:52]
  wire [11:0] _T_120; // @[Cat.scala 29:58]
  wire [11:0] _T_121; // @[Shift.scala 64:27]
  wire [1:0] _T_122; // @[Shift.scala 66:70]
  wire  _T_123; // @[Shift.scala 12:21]
  wire [9:0] _T_124; // @[Shift.scala 64:52]
  wire [11:0] _T_126; // @[Cat.scala 29:58]
  wire [11:0] _T_127; // @[Shift.scala 64:27]
  wire  _T_128; // @[Shift.scala 66:70]
  wire [10:0] _T_130; // @[Shift.scala 64:52]
  wire [11:0] _T_131; // @[Cat.scala 29:58]
  wire [11:0] _T_132; // @[Shift.scala 64:27]
  wire [11:0] _T_133; // @[Shift.scala 16:10]
  wire  _T_134; // @[convert.scala 23:34]
  wire [10:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_136; // @[convert.scala 25:26]
  wire [3:0] _T_138; // @[convert.scala 25:42]
  wire  _T_141; // @[convert.scala 26:67]
  wire  _T_142; // @[convert.scala 26:51]
  wire [5:0] _T_143; // @[Cat.scala 29:58]
  wire [13:0] _T_145; // @[convert.scala 29:56]
  wire  _T_146; // @[convert.scala 29:60]
  wire  _T_147; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_150; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_159; // @[convert.scala 18:24]
  wire  _T_160; // @[convert.scala 18:40]
  wire  _T_161; // @[convert.scala 18:36]
  wire [12:0] _T_162; // @[convert.scala 19:24]
  wire [12:0] _T_163; // @[convert.scala 19:43]
  wire [12:0] _T_164; // @[convert.scala 19:39]
  wire [7:0] _T_165; // @[LZD.scala 43:32]
  wire [3:0] _T_166; // @[LZD.scala 43:32]
  wire [1:0] _T_167; // @[LZD.scala 43:32]
  wire  _T_168; // @[LZD.scala 39:14]
  wire  _T_169; // @[LZD.scala 39:21]
  wire  _T_170; // @[LZD.scala 39:30]
  wire  _T_171; // @[LZD.scala 39:27]
  wire  _T_172; // @[LZD.scala 39:25]
  wire [1:0] _T_173; // @[Cat.scala 29:58]
  wire [1:0] _T_174; // @[LZD.scala 44:32]
  wire  _T_175; // @[LZD.scala 39:14]
  wire  _T_176; // @[LZD.scala 39:21]
  wire  _T_177; // @[LZD.scala 39:30]
  wire  _T_178; // @[LZD.scala 39:27]
  wire  _T_179; // @[LZD.scala 39:25]
  wire [1:0] _T_180; // @[Cat.scala 29:58]
  wire  _T_181; // @[Shift.scala 12:21]
  wire  _T_182; // @[Shift.scala 12:21]
  wire  _T_183; // @[LZD.scala 49:16]
  wire  _T_184; // @[LZD.scala 49:27]
  wire  _T_185; // @[LZD.scala 49:25]
  wire  _T_186; // @[LZD.scala 49:47]
  wire  _T_187; // @[LZD.scala 49:59]
  wire  _T_188; // @[LZD.scala 49:35]
  wire [2:0] _T_190; // @[Cat.scala 29:58]
  wire [3:0] _T_191; // @[LZD.scala 44:32]
  wire [1:0] _T_192; // @[LZD.scala 43:32]
  wire  _T_193; // @[LZD.scala 39:14]
  wire  _T_194; // @[LZD.scala 39:21]
  wire  _T_195; // @[LZD.scala 39:30]
  wire  _T_196; // @[LZD.scala 39:27]
  wire  _T_197; // @[LZD.scala 39:25]
  wire [1:0] _T_198; // @[Cat.scala 29:58]
  wire [1:0] _T_199; // @[LZD.scala 44:32]
  wire  _T_200; // @[LZD.scala 39:14]
  wire  _T_201; // @[LZD.scala 39:21]
  wire  _T_202; // @[LZD.scala 39:30]
  wire  _T_203; // @[LZD.scala 39:27]
  wire  _T_204; // @[LZD.scala 39:25]
  wire [1:0] _T_205; // @[Cat.scala 29:58]
  wire  _T_206; // @[Shift.scala 12:21]
  wire  _T_207; // @[Shift.scala 12:21]
  wire  _T_208; // @[LZD.scala 49:16]
  wire  _T_209; // @[LZD.scala 49:27]
  wire  _T_210; // @[LZD.scala 49:25]
  wire  _T_211; // @[LZD.scala 49:47]
  wire  _T_212; // @[LZD.scala 49:59]
  wire  _T_213; // @[LZD.scala 49:35]
  wire [2:0] _T_215; // @[Cat.scala 29:58]
  wire  _T_216; // @[Shift.scala 12:21]
  wire  _T_217; // @[Shift.scala 12:21]
  wire  _T_218; // @[LZD.scala 49:16]
  wire  _T_219; // @[LZD.scala 49:27]
  wire  _T_220; // @[LZD.scala 49:25]
  wire [1:0] _T_221; // @[LZD.scala 49:47]
  wire [1:0] _T_222; // @[LZD.scala 49:59]
  wire [1:0] _T_223; // @[LZD.scala 49:35]
  wire [3:0] _T_225; // @[Cat.scala 29:58]
  wire [4:0] _T_226; // @[LZD.scala 44:32]
  wire [3:0] _T_227; // @[LZD.scala 43:32]
  wire [1:0] _T_228; // @[LZD.scala 43:32]
  wire  _T_229; // @[LZD.scala 39:14]
  wire  _T_230; // @[LZD.scala 39:21]
  wire  _T_231; // @[LZD.scala 39:30]
  wire  _T_232; // @[LZD.scala 39:27]
  wire  _T_233; // @[LZD.scala 39:25]
  wire [1:0] _T_234; // @[Cat.scala 29:58]
  wire [1:0] _T_235; // @[LZD.scala 44:32]
  wire  _T_236; // @[LZD.scala 39:14]
  wire  _T_237; // @[LZD.scala 39:21]
  wire  _T_238; // @[LZD.scala 39:30]
  wire  _T_239; // @[LZD.scala 39:27]
  wire  _T_240; // @[LZD.scala 39:25]
  wire [1:0] _T_241; // @[Cat.scala 29:58]
  wire  _T_242; // @[Shift.scala 12:21]
  wire  _T_243; // @[Shift.scala 12:21]
  wire  _T_244; // @[LZD.scala 49:16]
  wire  _T_245; // @[LZD.scala 49:27]
  wire  _T_246; // @[LZD.scala 49:25]
  wire  _T_247; // @[LZD.scala 49:47]
  wire  _T_248; // @[LZD.scala 49:59]
  wire  _T_249; // @[LZD.scala 49:35]
  wire [2:0] _T_251; // @[Cat.scala 29:58]
  wire  _T_252; // @[LZD.scala 44:32]
  wire  _T_254; // @[Shift.scala 12:21]
  wire [1:0] _T_256; // @[Cat.scala 29:58]
  wire [1:0] _T_257; // @[LZD.scala 55:32]
  wire [1:0] _T_258; // @[LZD.scala 55:20]
  wire [2:0] _T_259; // @[Cat.scala 29:58]
  wire  _T_260; // @[Shift.scala 12:21]
  wire [2:0] _T_262; // @[LZD.scala 55:32]
  wire [2:0] _T_263; // @[LZD.scala 55:20]
  wire [3:0] _T_264; // @[Cat.scala 29:58]
  wire [3:0] _T_265; // @[convert.scala 21:22]
  wire [11:0] _T_266; // @[convert.scala 22:36]
  wire  _T_267; // @[Shift.scala 16:24]
  wire  _T_269; // @[Shift.scala 12:21]
  wire [3:0] _T_270; // @[Shift.scala 64:52]
  wire [11:0] _T_272; // @[Cat.scala 29:58]
  wire [11:0] _T_273; // @[Shift.scala 64:27]
  wire [2:0] _T_274; // @[Shift.scala 66:70]
  wire  _T_275; // @[Shift.scala 12:21]
  wire [7:0] _T_276; // @[Shift.scala 64:52]
  wire [11:0] _T_278; // @[Cat.scala 29:58]
  wire [11:0] _T_279; // @[Shift.scala 64:27]
  wire [1:0] _T_280; // @[Shift.scala 66:70]
  wire  _T_281; // @[Shift.scala 12:21]
  wire [9:0] _T_282; // @[Shift.scala 64:52]
  wire [11:0] _T_284; // @[Cat.scala 29:58]
  wire [11:0] _T_285; // @[Shift.scala 64:27]
  wire  _T_286; // @[Shift.scala 66:70]
  wire [10:0] _T_288; // @[Shift.scala 64:52]
  wire [11:0] _T_289; // @[Cat.scala 29:58]
  wire [11:0] _T_290; // @[Shift.scala 64:27]
  wire [11:0] _T_291; // @[Shift.scala 16:10]
  wire  _T_292; // @[convert.scala 23:34]
  wire [10:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_294; // @[convert.scala 25:26]
  wire [3:0] _T_296; // @[convert.scala 25:42]
  wire  _T_299; // @[convert.scala 26:67]
  wire  _T_300; // @[convert.scala 26:51]
  wire [5:0] _T_301; // @[Cat.scala 29:58]
  wire [13:0] _T_303; // @[convert.scala 29:56]
  wire  _T_304; // @[convert.scala 29:60]
  wire  _T_305; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_308; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  aGTb; // @[PositAdder.scala 24:32]
  wire  greaterSign; // @[PositAdder.scala 25:24]
  wire  smallerSign; // @[PositAdder.scala 26:24]
  wire [5:0] greaterExp; // @[PositAdder.scala 27:24]
  wire [5:0] smallerExp; // @[PositAdder.scala 28:24]
  wire [10:0] greaterFrac; // @[PositAdder.scala 29:24]
  wire [10:0] smallerFrac; // @[PositAdder.scala 30:24]
  wire [5:0] _T_317; // @[PositAdder.scala 31:32]
  wire [5:0] scale_diff; // @[PositAdder.scala 31:32]
  wire  _T_318; // @[PositAdder.scala 32:38]
  wire [12:0] greaterSig; // @[Cat.scala 29:58]
  wire  _T_320; // @[PositAdder.scala 33:38]
  wire [15:0] _T_323; // @[Cat.scala 29:58]
  wire [5:0] _T_324; // @[PositAdder.scala 34:68]
  wire  _T_325; // @[Shift.scala 39:24]
  wire [3:0] _T_326; // @[Shift.scala 40:44]
  wire [7:0] _T_327; // @[Shift.scala 90:30]
  wire [7:0] _T_328; // @[Shift.scala 90:48]
  wire  _T_329; // @[Shift.scala 90:57]
  wire [7:0] _GEN_0; // @[Shift.scala 90:39]
  wire [7:0] _T_330; // @[Shift.scala 90:39]
  wire  _T_331; // @[Shift.scala 12:21]
  wire  _T_332; // @[Shift.scala 12:21]
  wire [7:0] _T_334; // @[Bitwise.scala 71:12]
  wire [15:0] _T_335; // @[Cat.scala 29:58]
  wire [15:0] _T_336; // @[Shift.scala 91:22]
  wire [2:0] _T_337; // @[Shift.scala 92:77]
  wire [11:0] _T_338; // @[Shift.scala 90:30]
  wire [3:0] _T_339; // @[Shift.scala 90:48]
  wire  _T_340; // @[Shift.scala 90:57]
  wire [11:0] _GEN_1; // @[Shift.scala 90:39]
  wire [11:0] _T_341; // @[Shift.scala 90:39]
  wire  _T_342; // @[Shift.scala 12:21]
  wire  _T_343; // @[Shift.scala 12:21]
  wire [3:0] _T_345; // @[Bitwise.scala 71:12]
  wire [15:0] _T_346; // @[Cat.scala 29:58]
  wire [15:0] _T_347; // @[Shift.scala 91:22]
  wire [1:0] _T_348; // @[Shift.scala 92:77]
  wire [13:0] _T_349; // @[Shift.scala 90:30]
  wire [1:0] _T_350; // @[Shift.scala 90:48]
  wire  _T_351; // @[Shift.scala 90:57]
  wire [13:0] _GEN_2; // @[Shift.scala 90:39]
  wire [13:0] _T_352; // @[Shift.scala 90:39]
  wire  _T_353; // @[Shift.scala 12:21]
  wire  _T_354; // @[Shift.scala 12:21]
  wire [1:0] _T_356; // @[Bitwise.scala 71:12]
  wire [15:0] _T_357; // @[Cat.scala 29:58]
  wire [15:0] _T_358; // @[Shift.scala 91:22]
  wire  _T_359; // @[Shift.scala 92:77]
  wire [14:0] _T_360; // @[Shift.scala 90:30]
  wire  _T_361; // @[Shift.scala 90:48]
  wire [14:0] _GEN_3; // @[Shift.scala 90:39]
  wire [14:0] _T_363; // @[Shift.scala 90:39]
  wire  _T_365; // @[Shift.scala 12:21]
  wire [15:0] _T_366; // @[Cat.scala 29:58]
  wire [15:0] _T_367; // @[Shift.scala 91:22]
  wire [15:0] _T_370; // @[Bitwise.scala 71:12]
  wire [15:0] smallerSig; // @[Shift.scala 39:10]
  wire [12:0] _T_371; // @[PositAdder.scala 35:45]
  wire [13:0] rawSumSig; // @[PositAdder.scala 35:32]
  wire  _T_372; // @[PositAdder.scala 36:31]
  wire  _T_373; // @[PositAdder.scala 36:59]
  wire  sumSign; // @[PositAdder.scala 36:43]
  wire [12:0] _T_374; // @[PositAdder.scala 37:48]
  wire [2:0] _T_375; // @[PositAdder.scala 37:63]
  wire [16:0] signSumSig; // @[Cat.scala 29:58]
  wire [15:0] _T_377; // @[PositAdder.scala 39:31]
  wire [15:0] _T_378; // @[PositAdder.scala 39:66]
  wire [15:0] sumXor; // @[PositAdder.scala 39:49]
  wire [7:0] _T_379; // @[LZD.scala 43:32]
  wire [3:0] _T_380; // @[LZD.scala 43:32]
  wire [1:0] _T_381; // @[LZD.scala 43:32]
  wire  _T_382; // @[LZD.scala 39:14]
  wire  _T_383; // @[LZD.scala 39:21]
  wire  _T_384; // @[LZD.scala 39:30]
  wire  _T_385; // @[LZD.scala 39:27]
  wire  _T_386; // @[LZD.scala 39:25]
  wire [1:0] _T_387; // @[Cat.scala 29:58]
  wire [1:0] _T_388; // @[LZD.scala 44:32]
  wire  _T_389; // @[LZD.scala 39:14]
  wire  _T_390; // @[LZD.scala 39:21]
  wire  _T_391; // @[LZD.scala 39:30]
  wire  _T_392; // @[LZD.scala 39:27]
  wire  _T_393; // @[LZD.scala 39:25]
  wire [1:0] _T_394; // @[Cat.scala 29:58]
  wire  _T_395; // @[Shift.scala 12:21]
  wire  _T_396; // @[Shift.scala 12:21]
  wire  _T_397; // @[LZD.scala 49:16]
  wire  _T_398; // @[LZD.scala 49:27]
  wire  _T_399; // @[LZD.scala 49:25]
  wire  _T_400; // @[LZD.scala 49:47]
  wire  _T_401; // @[LZD.scala 49:59]
  wire  _T_402; // @[LZD.scala 49:35]
  wire [2:0] _T_404; // @[Cat.scala 29:58]
  wire [3:0] _T_405; // @[LZD.scala 44:32]
  wire [1:0] _T_406; // @[LZD.scala 43:32]
  wire  _T_407; // @[LZD.scala 39:14]
  wire  _T_408; // @[LZD.scala 39:21]
  wire  _T_409; // @[LZD.scala 39:30]
  wire  _T_410; // @[LZD.scala 39:27]
  wire  _T_411; // @[LZD.scala 39:25]
  wire [1:0] _T_412; // @[Cat.scala 29:58]
  wire [1:0] _T_413; // @[LZD.scala 44:32]
  wire  _T_414; // @[LZD.scala 39:14]
  wire  _T_415; // @[LZD.scala 39:21]
  wire  _T_416; // @[LZD.scala 39:30]
  wire  _T_417; // @[LZD.scala 39:27]
  wire  _T_418; // @[LZD.scala 39:25]
  wire [1:0] _T_419; // @[Cat.scala 29:58]
  wire  _T_420; // @[Shift.scala 12:21]
  wire  _T_421; // @[Shift.scala 12:21]
  wire  _T_422; // @[LZD.scala 49:16]
  wire  _T_423; // @[LZD.scala 49:27]
  wire  _T_424; // @[LZD.scala 49:25]
  wire  _T_425; // @[LZD.scala 49:47]
  wire  _T_426; // @[LZD.scala 49:59]
  wire  _T_427; // @[LZD.scala 49:35]
  wire [2:0] _T_429; // @[Cat.scala 29:58]
  wire  _T_430; // @[Shift.scala 12:21]
  wire  _T_431; // @[Shift.scala 12:21]
  wire  _T_432; // @[LZD.scala 49:16]
  wire  _T_433; // @[LZD.scala 49:27]
  wire  _T_434; // @[LZD.scala 49:25]
  wire [1:0] _T_435; // @[LZD.scala 49:47]
  wire [1:0] _T_436; // @[LZD.scala 49:59]
  wire [1:0] _T_437; // @[LZD.scala 49:35]
  wire [3:0] _T_439; // @[Cat.scala 29:58]
  wire [7:0] _T_440; // @[LZD.scala 44:32]
  wire [3:0] _T_441; // @[LZD.scala 43:32]
  wire [1:0] _T_442; // @[LZD.scala 43:32]
  wire  _T_443; // @[LZD.scala 39:14]
  wire  _T_444; // @[LZD.scala 39:21]
  wire  _T_445; // @[LZD.scala 39:30]
  wire  _T_446; // @[LZD.scala 39:27]
  wire  _T_447; // @[LZD.scala 39:25]
  wire [1:0] _T_448; // @[Cat.scala 29:58]
  wire [1:0] _T_449; // @[LZD.scala 44:32]
  wire  _T_450; // @[LZD.scala 39:14]
  wire  _T_451; // @[LZD.scala 39:21]
  wire  _T_452; // @[LZD.scala 39:30]
  wire  _T_453; // @[LZD.scala 39:27]
  wire  _T_454; // @[LZD.scala 39:25]
  wire [1:0] _T_455; // @[Cat.scala 29:58]
  wire  _T_456; // @[Shift.scala 12:21]
  wire  _T_457; // @[Shift.scala 12:21]
  wire  _T_458; // @[LZD.scala 49:16]
  wire  _T_459; // @[LZD.scala 49:27]
  wire  _T_460; // @[LZD.scala 49:25]
  wire  _T_461; // @[LZD.scala 49:47]
  wire  _T_462; // @[LZD.scala 49:59]
  wire  _T_463; // @[LZD.scala 49:35]
  wire [2:0] _T_465; // @[Cat.scala 29:58]
  wire [3:0] _T_466; // @[LZD.scala 44:32]
  wire [1:0] _T_467; // @[LZD.scala 43:32]
  wire  _T_468; // @[LZD.scala 39:14]
  wire  _T_469; // @[LZD.scala 39:21]
  wire  _T_470; // @[LZD.scala 39:30]
  wire  _T_471; // @[LZD.scala 39:27]
  wire  _T_472; // @[LZD.scala 39:25]
  wire [1:0] _T_473; // @[Cat.scala 29:58]
  wire [1:0] _T_474; // @[LZD.scala 44:32]
  wire  _T_475; // @[LZD.scala 39:14]
  wire  _T_476; // @[LZD.scala 39:21]
  wire  _T_477; // @[LZD.scala 39:30]
  wire  _T_478; // @[LZD.scala 39:27]
  wire  _T_479; // @[LZD.scala 39:25]
  wire [1:0] _T_480; // @[Cat.scala 29:58]
  wire  _T_481; // @[Shift.scala 12:21]
  wire  _T_482; // @[Shift.scala 12:21]
  wire  _T_483; // @[LZD.scala 49:16]
  wire  _T_484; // @[LZD.scala 49:27]
  wire  _T_485; // @[LZD.scala 49:25]
  wire  _T_486; // @[LZD.scala 49:47]
  wire  _T_487; // @[LZD.scala 49:59]
  wire  _T_488; // @[LZD.scala 49:35]
  wire [2:0] _T_490; // @[Cat.scala 29:58]
  wire  _T_491; // @[Shift.scala 12:21]
  wire  _T_492; // @[Shift.scala 12:21]
  wire  _T_493; // @[LZD.scala 49:16]
  wire  _T_494; // @[LZD.scala 49:27]
  wire  _T_495; // @[LZD.scala 49:25]
  wire [1:0] _T_496; // @[LZD.scala 49:47]
  wire [1:0] _T_497; // @[LZD.scala 49:59]
  wire [1:0] _T_498; // @[LZD.scala 49:35]
  wire [3:0] _T_500; // @[Cat.scala 29:58]
  wire  _T_501; // @[Shift.scala 12:21]
  wire  _T_502; // @[Shift.scala 12:21]
  wire  _T_503; // @[LZD.scala 49:16]
  wire  _T_504; // @[LZD.scala 49:27]
  wire  _T_505; // @[LZD.scala 49:25]
  wire [2:0] _T_506; // @[LZD.scala 49:47]
  wire [2:0] _T_507; // @[LZD.scala 49:59]
  wire [2:0] _T_508; // @[LZD.scala 49:35]
  wire [4:0] sumLZD; // @[Cat.scala 29:58]
  wire [5:0] _T_510; // @[Cat.scala 29:58]
  wire [5:0] _T_511; // @[PositAdder.scala 41:38]
  wire [5:0] _T_513; // @[PositAdder.scala 41:45]
  wire [5:0] scaleBias; // @[PositAdder.scala 41:45]
  wire [6:0] sumScale; // @[PositAdder.scala 42:32]
  wire  overflow; // @[PositAdder.scala 43:30]
  wire [4:0] normalShift; // @[PositAdder.scala 44:22]
  wire [14:0] _T_514; // @[PositAdder.scala 45:36]
  wire  _T_515; // @[Shift.scala 16:24]
  wire [3:0] _T_516; // @[Shift.scala 17:37]
  wire  _T_517; // @[Shift.scala 12:21]
  wire [6:0] _T_518; // @[Shift.scala 64:52]
  wire [14:0] _T_520; // @[Cat.scala 29:58]
  wire [14:0] _T_521; // @[Shift.scala 64:27]
  wire [2:0] _T_522; // @[Shift.scala 66:70]
  wire  _T_523; // @[Shift.scala 12:21]
  wire [10:0] _T_524; // @[Shift.scala 64:52]
  wire [14:0] _T_526; // @[Cat.scala 29:58]
  wire [14:0] _T_527; // @[Shift.scala 64:27]
  wire [1:0] _T_528; // @[Shift.scala 66:70]
  wire  _T_529; // @[Shift.scala 12:21]
  wire [12:0] _T_530; // @[Shift.scala 64:52]
  wire [14:0] _T_532; // @[Cat.scala 29:58]
  wire [14:0] _T_533; // @[Shift.scala 64:27]
  wire  _T_534; // @[Shift.scala 66:70]
  wire [13:0] _T_536; // @[Shift.scala 64:52]
  wire [14:0] _T_537; // @[Cat.scala 29:58]
  wire [14:0] _T_538; // @[Shift.scala 64:27]
  wire [14:0] shiftSig; // @[Shift.scala 16:10]
  wire [6:0] _T_539; // @[PositAdder.scala 50:24]
  wire [10:0] decS_fraction; // @[PositAdder.scala 51:34]
  wire  decS_isNaR; // @[PositAdder.scala 52:32]
  wire  _T_542; // @[PositAdder.scala 53:33]
  wire  _T_543; // @[PositAdder.scala 53:21]
  wire  _T_544; // @[PositAdder.scala 53:52]
  wire  decS_isZero; // @[PositAdder.scala 53:37]
  wire [1:0] _T_546; // @[PositAdder.scala 54:33]
  wire  _T_547; // @[PositAdder.scala 54:49]
  wire  _T_548; // @[PositAdder.scala 54:63]
  wire  _T_549; // @[PositAdder.scala 54:53]
  wire [5:0] _GEN_4; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  wire [5:0] decS_scale; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  wire  _T_552; // @[convert.scala 46:61]
  wire  _T_553; // @[convert.scala 46:52]
  wire  _T_555; // @[convert.scala 46:42]
  wire [4:0] _T_556; // @[convert.scala 48:34]
  wire  _T_557; // @[convert.scala 49:36]
  wire [4:0] _T_559; // @[convert.scala 50:36]
  wire [4:0] _T_560; // @[convert.scala 50:36]
  wire [4:0] _T_561; // @[convert.scala 50:28]
  wire  _T_562; // @[convert.scala 51:31]
  wire  _T_563; // @[convert.scala 52:43]
  wire [16:0] _T_567; // @[Cat.scala 29:58]
  wire [4:0] _T_568; // @[Shift.scala 39:17]
  wire  _T_569; // @[Shift.scala 39:24]
  wire  _T_571; // @[Shift.scala 90:30]
  wire [15:0] _T_572; // @[Shift.scala 90:48]
  wire  _T_573; // @[Shift.scala 90:57]
  wire  _T_574; // @[Shift.scala 90:39]
  wire  _T_575; // @[Shift.scala 12:21]
  wire  _T_576; // @[Shift.scala 12:21]
  wire [15:0] _T_578; // @[Bitwise.scala 71:12]
  wire [16:0] _T_579; // @[Cat.scala 29:58]
  wire [16:0] _T_580; // @[Shift.scala 91:22]
  wire [3:0] _T_581; // @[Shift.scala 92:77]
  wire [8:0] _T_582; // @[Shift.scala 90:30]
  wire [7:0] _T_583; // @[Shift.scala 90:48]
  wire  _T_584; // @[Shift.scala 90:57]
  wire [8:0] _GEN_5; // @[Shift.scala 90:39]
  wire [8:0] _T_585; // @[Shift.scala 90:39]
  wire  _T_586; // @[Shift.scala 12:21]
  wire  _T_587; // @[Shift.scala 12:21]
  wire [7:0] _T_589; // @[Bitwise.scala 71:12]
  wire [16:0] _T_590; // @[Cat.scala 29:58]
  wire [16:0] _T_591; // @[Shift.scala 91:22]
  wire [2:0] _T_592; // @[Shift.scala 92:77]
  wire [12:0] _T_593; // @[Shift.scala 90:30]
  wire [3:0] _T_594; // @[Shift.scala 90:48]
  wire  _T_595; // @[Shift.scala 90:57]
  wire [12:0] _GEN_6; // @[Shift.scala 90:39]
  wire [12:0] _T_596; // @[Shift.scala 90:39]
  wire  _T_597; // @[Shift.scala 12:21]
  wire  _T_598; // @[Shift.scala 12:21]
  wire [3:0] _T_600; // @[Bitwise.scala 71:12]
  wire [16:0] _T_601; // @[Cat.scala 29:58]
  wire [16:0] _T_602; // @[Shift.scala 91:22]
  wire [1:0] _T_603; // @[Shift.scala 92:77]
  wire [14:0] _T_604; // @[Shift.scala 90:30]
  wire [1:0] _T_605; // @[Shift.scala 90:48]
  wire  _T_606; // @[Shift.scala 90:57]
  wire [14:0] _GEN_7; // @[Shift.scala 90:39]
  wire [14:0] _T_607; // @[Shift.scala 90:39]
  wire  _T_608; // @[Shift.scala 12:21]
  wire  _T_609; // @[Shift.scala 12:21]
  wire [1:0] _T_611; // @[Bitwise.scala 71:12]
  wire [16:0] _T_612; // @[Cat.scala 29:58]
  wire [16:0] _T_613; // @[Shift.scala 91:22]
  wire  _T_614; // @[Shift.scala 92:77]
  wire [15:0] _T_615; // @[Shift.scala 90:30]
  wire  _T_616; // @[Shift.scala 90:48]
  wire [15:0] _GEN_8; // @[Shift.scala 90:39]
  wire [15:0] _T_618; // @[Shift.scala 90:39]
  wire  _T_620; // @[Shift.scala 12:21]
  wire [16:0] _T_621; // @[Cat.scala 29:58]
  wire [16:0] _T_622; // @[Shift.scala 91:22]
  wire [16:0] _T_625; // @[Bitwise.scala 71:12]
  wire [16:0] _T_626; // @[Shift.scala 39:10]
  wire  _T_627; // @[convert.scala 55:31]
  wire  _T_628; // @[convert.scala 56:31]
  wire  _T_629; // @[convert.scala 57:31]
  wire  _T_630; // @[convert.scala 58:31]
  wire [13:0] _T_631; // @[convert.scala 59:69]
  wire  _T_632; // @[convert.scala 59:81]
  wire  _T_633; // @[convert.scala 59:50]
  wire  _T_635; // @[convert.scala 60:81]
  wire  _T_636; // @[convert.scala 61:44]
  wire  _T_637; // @[convert.scala 61:52]
  wire  _T_638; // @[convert.scala 61:36]
  wire  _T_639; // @[convert.scala 62:63]
  wire  _T_640; // @[convert.scala 62:103]
  wire  _T_641; // @[convert.scala 62:60]
  wire [13:0] _GEN_9; // @[convert.scala 63:56]
  wire [13:0] _T_644; // @[convert.scala 63:56]
  wire [14:0] _T_645; // @[Cat.scala 29:58]
  wire [14:0] _T_647; // @[Mux.scala 87:16]
  assign _T_1 = io_A[14]; // @[convert.scala 18:24]
  assign _T_2 = io_A[13]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[13:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[12:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[12:5]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[4:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68[4:1]; // @[LZD.scala 43:32]
  assign _T_70 = _T_69[3:2]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70 != 2'h0; // @[LZD.scala 39:14]
  assign _T_72 = _T_70[1]; // @[LZD.scala 39:21]
  assign _T_73 = _T_70[0]; // @[LZD.scala 39:30]
  assign _T_74 = ~ _T_73; // @[LZD.scala 39:27]
  assign _T_75 = _T_72 | _T_74; // @[LZD.scala 39:25]
  assign _T_76 = {_T_71,_T_75}; // @[Cat.scala 29:58]
  assign _T_77 = _T_69[1:0]; // @[LZD.scala 44:32]
  assign _T_78 = _T_77 != 2'h0; // @[LZD.scala 39:14]
  assign _T_79 = _T_77[1]; // @[LZD.scala 39:21]
  assign _T_80 = _T_77[0]; // @[LZD.scala 39:30]
  assign _T_81 = ~ _T_80; // @[LZD.scala 39:27]
  assign _T_82 = _T_79 | _T_81; // @[LZD.scala 39:25]
  assign _T_83 = {_T_78,_T_82}; // @[Cat.scala 29:58]
  assign _T_84 = _T_76[1]; // @[Shift.scala 12:21]
  assign _T_85 = _T_83[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84 | _T_85; // @[LZD.scala 49:16]
  assign _T_87 = ~ _T_85; // @[LZD.scala 49:27]
  assign _T_88 = _T_84 | _T_87; // @[LZD.scala 49:25]
  assign _T_89 = _T_76[0:0]; // @[LZD.scala 49:47]
  assign _T_90 = _T_83[0:0]; // @[LZD.scala 49:59]
  assign _T_91 = _T_84 ? _T_89 : _T_90; // @[LZD.scala 49:35]
  assign _T_93 = {_T_86,_T_88,_T_91}; // @[Cat.scala 29:58]
  assign _T_94 = _T_68[0:0]; // @[LZD.scala 44:32]
  assign _T_96 = _T_93[2]; // @[Shift.scala 12:21]
  assign _T_98 = {1'h1,_T_94}; // @[Cat.scala 29:58]
  assign _T_99 = _T_93[1:0]; // @[LZD.scala 55:32]
  assign _T_100 = _T_96 ? _T_99 : _T_98; // @[LZD.scala 55:20]
  assign _T_101 = {_T_96,_T_100}; // @[Cat.scala 29:58]
  assign _T_102 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_104 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_105 = _T_102 ? _T_104 : _T_101; // @[LZD.scala 55:20]
  assign _T_106 = {_T_102,_T_105}; // @[Cat.scala 29:58]
  assign _T_107 = ~ _T_106; // @[convert.scala 21:22]
  assign _T_108 = io_A[11:0]; // @[convert.scala 22:36]
  assign _T_109 = _T_107 < 4'hc; // @[Shift.scala 16:24]
  assign _T_111 = _T_107[3]; // @[Shift.scala 12:21]
  assign _T_112 = _T_108[3:0]; // @[Shift.scala 64:52]
  assign _T_114 = {_T_112,8'h0}; // @[Cat.scala 29:58]
  assign _T_115 = _T_111 ? _T_114 : _T_108; // @[Shift.scala 64:27]
  assign _T_116 = _T_107[2:0]; // @[Shift.scala 66:70]
  assign _T_117 = _T_116[2]; // @[Shift.scala 12:21]
  assign _T_118 = _T_115[7:0]; // @[Shift.scala 64:52]
  assign _T_120 = {_T_118,4'h0}; // @[Cat.scala 29:58]
  assign _T_121 = _T_117 ? _T_120 : _T_115; // @[Shift.scala 64:27]
  assign _T_122 = _T_116[1:0]; // @[Shift.scala 66:70]
  assign _T_123 = _T_122[1]; // @[Shift.scala 12:21]
  assign _T_124 = _T_121[9:0]; // @[Shift.scala 64:52]
  assign _T_126 = {_T_124,2'h0}; // @[Cat.scala 29:58]
  assign _T_127 = _T_123 ? _T_126 : _T_121; // @[Shift.scala 64:27]
  assign _T_128 = _T_122[0:0]; // @[Shift.scala 66:70]
  assign _T_130 = _T_127[10:0]; // @[Shift.scala 64:52]
  assign _T_131 = {_T_130,1'h0}; // @[Cat.scala 29:58]
  assign _T_132 = _T_128 ? _T_131 : _T_127; // @[Shift.scala 64:27]
  assign _T_133 = _T_109 ? _T_132 : 12'h0; // @[Shift.scala 16:10]
  assign _T_134 = _T_133[11:11]; // @[convert.scala 23:34]
  assign decA_fraction = _T_133[10:0]; // @[convert.scala 24:34]
  assign _T_136 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_138 = _T_3 ? _T_107 : _T_106; // @[convert.scala 25:42]
  assign _T_141 = ~ _T_134; // @[convert.scala 26:67]
  assign _T_142 = _T_1 ? _T_141 : _T_134; // @[convert.scala 26:51]
  assign _T_143 = {_T_136,_T_138,_T_142}; // @[Cat.scala 29:58]
  assign _T_145 = io_A[13:0]; // @[convert.scala 29:56]
  assign _T_146 = _T_145 != 14'h0; // @[convert.scala 29:60]
  assign _T_147 = ~ _T_146; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_147; // @[convert.scala 29:39]
  assign _T_150 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_150 & _T_147; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_143); // @[convert.scala 32:24]
  assign _T_159 = io_B[14]; // @[convert.scala 18:24]
  assign _T_160 = io_B[13]; // @[convert.scala 18:40]
  assign _T_161 = _T_159 ^ _T_160; // @[convert.scala 18:36]
  assign _T_162 = io_B[13:1]; // @[convert.scala 19:24]
  assign _T_163 = io_B[12:0]; // @[convert.scala 19:43]
  assign _T_164 = _T_162 ^ _T_163; // @[convert.scala 19:39]
  assign _T_165 = _T_164[12:5]; // @[LZD.scala 43:32]
  assign _T_166 = _T_165[7:4]; // @[LZD.scala 43:32]
  assign _T_167 = _T_166[3:2]; // @[LZD.scala 43:32]
  assign _T_168 = _T_167 != 2'h0; // @[LZD.scala 39:14]
  assign _T_169 = _T_167[1]; // @[LZD.scala 39:21]
  assign _T_170 = _T_167[0]; // @[LZD.scala 39:30]
  assign _T_171 = ~ _T_170; // @[LZD.scala 39:27]
  assign _T_172 = _T_169 | _T_171; // @[LZD.scala 39:25]
  assign _T_173 = {_T_168,_T_172}; // @[Cat.scala 29:58]
  assign _T_174 = _T_166[1:0]; // @[LZD.scala 44:32]
  assign _T_175 = _T_174 != 2'h0; // @[LZD.scala 39:14]
  assign _T_176 = _T_174[1]; // @[LZD.scala 39:21]
  assign _T_177 = _T_174[0]; // @[LZD.scala 39:30]
  assign _T_178 = ~ _T_177; // @[LZD.scala 39:27]
  assign _T_179 = _T_176 | _T_178; // @[LZD.scala 39:25]
  assign _T_180 = {_T_175,_T_179}; // @[Cat.scala 29:58]
  assign _T_181 = _T_173[1]; // @[Shift.scala 12:21]
  assign _T_182 = _T_180[1]; // @[Shift.scala 12:21]
  assign _T_183 = _T_181 | _T_182; // @[LZD.scala 49:16]
  assign _T_184 = ~ _T_182; // @[LZD.scala 49:27]
  assign _T_185 = _T_181 | _T_184; // @[LZD.scala 49:25]
  assign _T_186 = _T_173[0:0]; // @[LZD.scala 49:47]
  assign _T_187 = _T_180[0:0]; // @[LZD.scala 49:59]
  assign _T_188 = _T_181 ? _T_186 : _T_187; // @[LZD.scala 49:35]
  assign _T_190 = {_T_183,_T_185,_T_188}; // @[Cat.scala 29:58]
  assign _T_191 = _T_165[3:0]; // @[LZD.scala 44:32]
  assign _T_192 = _T_191[3:2]; // @[LZD.scala 43:32]
  assign _T_193 = _T_192 != 2'h0; // @[LZD.scala 39:14]
  assign _T_194 = _T_192[1]; // @[LZD.scala 39:21]
  assign _T_195 = _T_192[0]; // @[LZD.scala 39:30]
  assign _T_196 = ~ _T_195; // @[LZD.scala 39:27]
  assign _T_197 = _T_194 | _T_196; // @[LZD.scala 39:25]
  assign _T_198 = {_T_193,_T_197}; // @[Cat.scala 29:58]
  assign _T_199 = _T_191[1:0]; // @[LZD.scala 44:32]
  assign _T_200 = _T_199 != 2'h0; // @[LZD.scala 39:14]
  assign _T_201 = _T_199[1]; // @[LZD.scala 39:21]
  assign _T_202 = _T_199[0]; // @[LZD.scala 39:30]
  assign _T_203 = ~ _T_202; // @[LZD.scala 39:27]
  assign _T_204 = _T_201 | _T_203; // @[LZD.scala 39:25]
  assign _T_205 = {_T_200,_T_204}; // @[Cat.scala 29:58]
  assign _T_206 = _T_198[1]; // @[Shift.scala 12:21]
  assign _T_207 = _T_205[1]; // @[Shift.scala 12:21]
  assign _T_208 = _T_206 | _T_207; // @[LZD.scala 49:16]
  assign _T_209 = ~ _T_207; // @[LZD.scala 49:27]
  assign _T_210 = _T_206 | _T_209; // @[LZD.scala 49:25]
  assign _T_211 = _T_198[0:0]; // @[LZD.scala 49:47]
  assign _T_212 = _T_205[0:0]; // @[LZD.scala 49:59]
  assign _T_213 = _T_206 ? _T_211 : _T_212; // @[LZD.scala 49:35]
  assign _T_215 = {_T_208,_T_210,_T_213}; // @[Cat.scala 29:58]
  assign _T_216 = _T_190[2]; // @[Shift.scala 12:21]
  assign _T_217 = _T_215[2]; // @[Shift.scala 12:21]
  assign _T_218 = _T_216 | _T_217; // @[LZD.scala 49:16]
  assign _T_219 = ~ _T_217; // @[LZD.scala 49:27]
  assign _T_220 = _T_216 | _T_219; // @[LZD.scala 49:25]
  assign _T_221 = _T_190[1:0]; // @[LZD.scala 49:47]
  assign _T_222 = _T_215[1:0]; // @[LZD.scala 49:59]
  assign _T_223 = _T_216 ? _T_221 : _T_222; // @[LZD.scala 49:35]
  assign _T_225 = {_T_218,_T_220,_T_223}; // @[Cat.scala 29:58]
  assign _T_226 = _T_164[4:0]; // @[LZD.scala 44:32]
  assign _T_227 = _T_226[4:1]; // @[LZD.scala 43:32]
  assign _T_228 = _T_227[3:2]; // @[LZD.scala 43:32]
  assign _T_229 = _T_228 != 2'h0; // @[LZD.scala 39:14]
  assign _T_230 = _T_228[1]; // @[LZD.scala 39:21]
  assign _T_231 = _T_228[0]; // @[LZD.scala 39:30]
  assign _T_232 = ~ _T_231; // @[LZD.scala 39:27]
  assign _T_233 = _T_230 | _T_232; // @[LZD.scala 39:25]
  assign _T_234 = {_T_229,_T_233}; // @[Cat.scala 29:58]
  assign _T_235 = _T_227[1:0]; // @[LZD.scala 44:32]
  assign _T_236 = _T_235 != 2'h0; // @[LZD.scala 39:14]
  assign _T_237 = _T_235[1]; // @[LZD.scala 39:21]
  assign _T_238 = _T_235[0]; // @[LZD.scala 39:30]
  assign _T_239 = ~ _T_238; // @[LZD.scala 39:27]
  assign _T_240 = _T_237 | _T_239; // @[LZD.scala 39:25]
  assign _T_241 = {_T_236,_T_240}; // @[Cat.scala 29:58]
  assign _T_242 = _T_234[1]; // @[Shift.scala 12:21]
  assign _T_243 = _T_241[1]; // @[Shift.scala 12:21]
  assign _T_244 = _T_242 | _T_243; // @[LZD.scala 49:16]
  assign _T_245 = ~ _T_243; // @[LZD.scala 49:27]
  assign _T_246 = _T_242 | _T_245; // @[LZD.scala 49:25]
  assign _T_247 = _T_234[0:0]; // @[LZD.scala 49:47]
  assign _T_248 = _T_241[0:0]; // @[LZD.scala 49:59]
  assign _T_249 = _T_242 ? _T_247 : _T_248; // @[LZD.scala 49:35]
  assign _T_251 = {_T_244,_T_246,_T_249}; // @[Cat.scala 29:58]
  assign _T_252 = _T_226[0:0]; // @[LZD.scala 44:32]
  assign _T_254 = _T_251[2]; // @[Shift.scala 12:21]
  assign _T_256 = {1'h1,_T_252}; // @[Cat.scala 29:58]
  assign _T_257 = _T_251[1:0]; // @[LZD.scala 55:32]
  assign _T_258 = _T_254 ? _T_257 : _T_256; // @[LZD.scala 55:20]
  assign _T_259 = {_T_254,_T_258}; // @[Cat.scala 29:58]
  assign _T_260 = _T_225[3]; // @[Shift.scala 12:21]
  assign _T_262 = _T_225[2:0]; // @[LZD.scala 55:32]
  assign _T_263 = _T_260 ? _T_262 : _T_259; // @[LZD.scala 55:20]
  assign _T_264 = {_T_260,_T_263}; // @[Cat.scala 29:58]
  assign _T_265 = ~ _T_264; // @[convert.scala 21:22]
  assign _T_266 = io_B[11:0]; // @[convert.scala 22:36]
  assign _T_267 = _T_265 < 4'hc; // @[Shift.scala 16:24]
  assign _T_269 = _T_265[3]; // @[Shift.scala 12:21]
  assign _T_270 = _T_266[3:0]; // @[Shift.scala 64:52]
  assign _T_272 = {_T_270,8'h0}; // @[Cat.scala 29:58]
  assign _T_273 = _T_269 ? _T_272 : _T_266; // @[Shift.scala 64:27]
  assign _T_274 = _T_265[2:0]; // @[Shift.scala 66:70]
  assign _T_275 = _T_274[2]; // @[Shift.scala 12:21]
  assign _T_276 = _T_273[7:0]; // @[Shift.scala 64:52]
  assign _T_278 = {_T_276,4'h0}; // @[Cat.scala 29:58]
  assign _T_279 = _T_275 ? _T_278 : _T_273; // @[Shift.scala 64:27]
  assign _T_280 = _T_274[1:0]; // @[Shift.scala 66:70]
  assign _T_281 = _T_280[1]; // @[Shift.scala 12:21]
  assign _T_282 = _T_279[9:0]; // @[Shift.scala 64:52]
  assign _T_284 = {_T_282,2'h0}; // @[Cat.scala 29:58]
  assign _T_285 = _T_281 ? _T_284 : _T_279; // @[Shift.scala 64:27]
  assign _T_286 = _T_280[0:0]; // @[Shift.scala 66:70]
  assign _T_288 = _T_285[10:0]; // @[Shift.scala 64:52]
  assign _T_289 = {_T_288,1'h0}; // @[Cat.scala 29:58]
  assign _T_290 = _T_286 ? _T_289 : _T_285; // @[Shift.scala 64:27]
  assign _T_291 = _T_267 ? _T_290 : 12'h0; // @[Shift.scala 16:10]
  assign _T_292 = _T_291[11:11]; // @[convert.scala 23:34]
  assign decB_fraction = _T_291[10:0]; // @[convert.scala 24:34]
  assign _T_294 = _T_161 == 1'h0; // @[convert.scala 25:26]
  assign _T_296 = _T_161 ? _T_265 : _T_264; // @[convert.scala 25:42]
  assign _T_299 = ~ _T_292; // @[convert.scala 26:67]
  assign _T_300 = _T_159 ? _T_299 : _T_292; // @[convert.scala 26:51]
  assign _T_301 = {_T_294,_T_296,_T_300}; // @[Cat.scala 29:58]
  assign _T_303 = io_B[13:0]; // @[convert.scala 29:56]
  assign _T_304 = _T_303 != 14'h0; // @[convert.scala 29:60]
  assign _T_305 = ~ _T_304; // @[convert.scala 29:41]
  assign decB_isNaR = _T_159 & _T_305; // @[convert.scala 29:39]
  assign _T_308 = _T_159 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_308 & _T_305; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_301); // @[convert.scala 32:24]
  assign aGTb = $signed(decA_scale) > $signed(decB_scale); // @[PositAdder.scala 24:32]
  assign greaterSign = aGTb ? _T_1 : _T_159; // @[PositAdder.scala 25:24]
  assign smallerSign = aGTb ? _T_159 : _T_1; // @[PositAdder.scala 26:24]
  assign greaterExp = aGTb ? $signed(decA_scale) : $signed(decB_scale); // @[PositAdder.scala 27:24]
  assign smallerExp = aGTb ? $signed(decB_scale) : $signed(decA_scale); // @[PositAdder.scala 28:24]
  assign greaterFrac = aGTb ? decA_fraction : decB_fraction; // @[PositAdder.scala 29:24]
  assign smallerFrac = aGTb ? decB_fraction : decA_fraction; // @[PositAdder.scala 30:24]
  assign _T_317 = $signed(greaterExp) - $signed(smallerExp); // @[PositAdder.scala 31:32]
  assign scale_diff = $signed(_T_317); // @[PositAdder.scala 31:32]
  assign _T_318 = ~ greaterSign; // @[PositAdder.scala 32:38]
  assign greaterSig = {greaterSign,_T_318,greaterFrac}; // @[Cat.scala 29:58]
  assign _T_320 = ~ smallerSign; // @[PositAdder.scala 33:38]
  assign _T_323 = {smallerSign,_T_320,smallerFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_324 = $unsigned(scale_diff); // @[PositAdder.scala 34:68]
  assign _T_325 = _T_324 < 6'h10; // @[Shift.scala 39:24]
  assign _T_326 = _T_324[3:0]; // @[Shift.scala 40:44]
  assign _T_327 = _T_323[15:8]; // @[Shift.scala 90:30]
  assign _T_328 = _T_323[7:0]; // @[Shift.scala 90:48]
  assign _T_329 = _T_328 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_0 = {{7'd0}, _T_329}; // @[Shift.scala 90:39]
  assign _T_330 = _T_327 | _GEN_0; // @[Shift.scala 90:39]
  assign _T_331 = _T_326[3]; // @[Shift.scala 12:21]
  assign _T_332 = _T_323[15]; // @[Shift.scala 12:21]
  assign _T_334 = _T_332 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_335 = {_T_334,_T_330}; // @[Cat.scala 29:58]
  assign _T_336 = _T_331 ? _T_335 : _T_323; // @[Shift.scala 91:22]
  assign _T_337 = _T_326[2:0]; // @[Shift.scala 92:77]
  assign _T_338 = _T_336[15:4]; // @[Shift.scala 90:30]
  assign _T_339 = _T_336[3:0]; // @[Shift.scala 90:48]
  assign _T_340 = _T_339 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_1 = {{11'd0}, _T_340}; // @[Shift.scala 90:39]
  assign _T_341 = _T_338 | _GEN_1; // @[Shift.scala 90:39]
  assign _T_342 = _T_337[2]; // @[Shift.scala 12:21]
  assign _T_343 = _T_336[15]; // @[Shift.scala 12:21]
  assign _T_345 = _T_343 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_346 = {_T_345,_T_341}; // @[Cat.scala 29:58]
  assign _T_347 = _T_342 ? _T_346 : _T_336; // @[Shift.scala 91:22]
  assign _T_348 = _T_337[1:0]; // @[Shift.scala 92:77]
  assign _T_349 = _T_347[15:2]; // @[Shift.scala 90:30]
  assign _T_350 = _T_347[1:0]; // @[Shift.scala 90:48]
  assign _T_351 = _T_350 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{13'd0}, _T_351}; // @[Shift.scala 90:39]
  assign _T_352 = _T_349 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_353 = _T_348[1]; // @[Shift.scala 12:21]
  assign _T_354 = _T_347[15]; // @[Shift.scala 12:21]
  assign _T_356 = _T_354 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_357 = {_T_356,_T_352}; // @[Cat.scala 29:58]
  assign _T_358 = _T_353 ? _T_357 : _T_347; // @[Shift.scala 91:22]
  assign _T_359 = _T_348[0:0]; // @[Shift.scala 92:77]
  assign _T_360 = _T_358[15:1]; // @[Shift.scala 90:30]
  assign _T_361 = _T_358[0:0]; // @[Shift.scala 90:48]
  assign _GEN_3 = {{14'd0}, _T_361}; // @[Shift.scala 90:39]
  assign _T_363 = _T_360 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_365 = _T_358[15]; // @[Shift.scala 12:21]
  assign _T_366 = {_T_365,_T_363}; // @[Cat.scala 29:58]
  assign _T_367 = _T_359 ? _T_366 : _T_358; // @[Shift.scala 91:22]
  assign _T_370 = _T_332 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_325 ? _T_367 : _T_370; // @[Shift.scala 39:10]
  assign _T_371 = smallerSig[15:3]; // @[PositAdder.scala 35:45]
  assign rawSumSig = greaterSig + _T_371; // @[PositAdder.scala 35:32]
  assign _T_372 = _T_1 ^ _T_159; // @[PositAdder.scala 36:31]
  assign _T_373 = rawSumSig[13:13]; // @[PositAdder.scala 36:59]
  assign sumSign = _T_372 ^ _T_373; // @[PositAdder.scala 36:43]
  assign _T_374 = greaterSig + _T_371; // @[PositAdder.scala 37:48]
  assign _T_375 = smallerSig[2:0]; // @[PositAdder.scala 37:63]
  assign signSumSig = {sumSign,_T_374,_T_375}; // @[Cat.scala 29:58]
  assign _T_377 = signSumSig[16:1]; // @[PositAdder.scala 39:31]
  assign _T_378 = signSumSig[15:0]; // @[PositAdder.scala 39:66]
  assign sumXor = _T_377 ^ _T_378; // @[PositAdder.scala 39:49]
  assign _T_379 = sumXor[15:8]; // @[LZD.scala 43:32]
  assign _T_380 = _T_379[7:4]; // @[LZD.scala 43:32]
  assign _T_381 = _T_380[3:2]; // @[LZD.scala 43:32]
  assign _T_382 = _T_381 != 2'h0; // @[LZD.scala 39:14]
  assign _T_383 = _T_381[1]; // @[LZD.scala 39:21]
  assign _T_384 = _T_381[0]; // @[LZD.scala 39:30]
  assign _T_385 = ~ _T_384; // @[LZD.scala 39:27]
  assign _T_386 = _T_383 | _T_385; // @[LZD.scala 39:25]
  assign _T_387 = {_T_382,_T_386}; // @[Cat.scala 29:58]
  assign _T_388 = _T_380[1:0]; // @[LZD.scala 44:32]
  assign _T_389 = _T_388 != 2'h0; // @[LZD.scala 39:14]
  assign _T_390 = _T_388[1]; // @[LZD.scala 39:21]
  assign _T_391 = _T_388[0]; // @[LZD.scala 39:30]
  assign _T_392 = ~ _T_391; // @[LZD.scala 39:27]
  assign _T_393 = _T_390 | _T_392; // @[LZD.scala 39:25]
  assign _T_394 = {_T_389,_T_393}; // @[Cat.scala 29:58]
  assign _T_395 = _T_387[1]; // @[Shift.scala 12:21]
  assign _T_396 = _T_394[1]; // @[Shift.scala 12:21]
  assign _T_397 = _T_395 | _T_396; // @[LZD.scala 49:16]
  assign _T_398 = ~ _T_396; // @[LZD.scala 49:27]
  assign _T_399 = _T_395 | _T_398; // @[LZD.scala 49:25]
  assign _T_400 = _T_387[0:0]; // @[LZD.scala 49:47]
  assign _T_401 = _T_394[0:0]; // @[LZD.scala 49:59]
  assign _T_402 = _T_395 ? _T_400 : _T_401; // @[LZD.scala 49:35]
  assign _T_404 = {_T_397,_T_399,_T_402}; // @[Cat.scala 29:58]
  assign _T_405 = _T_379[3:0]; // @[LZD.scala 44:32]
  assign _T_406 = _T_405[3:2]; // @[LZD.scala 43:32]
  assign _T_407 = _T_406 != 2'h0; // @[LZD.scala 39:14]
  assign _T_408 = _T_406[1]; // @[LZD.scala 39:21]
  assign _T_409 = _T_406[0]; // @[LZD.scala 39:30]
  assign _T_410 = ~ _T_409; // @[LZD.scala 39:27]
  assign _T_411 = _T_408 | _T_410; // @[LZD.scala 39:25]
  assign _T_412 = {_T_407,_T_411}; // @[Cat.scala 29:58]
  assign _T_413 = _T_405[1:0]; // @[LZD.scala 44:32]
  assign _T_414 = _T_413 != 2'h0; // @[LZD.scala 39:14]
  assign _T_415 = _T_413[1]; // @[LZD.scala 39:21]
  assign _T_416 = _T_413[0]; // @[LZD.scala 39:30]
  assign _T_417 = ~ _T_416; // @[LZD.scala 39:27]
  assign _T_418 = _T_415 | _T_417; // @[LZD.scala 39:25]
  assign _T_419 = {_T_414,_T_418}; // @[Cat.scala 29:58]
  assign _T_420 = _T_412[1]; // @[Shift.scala 12:21]
  assign _T_421 = _T_419[1]; // @[Shift.scala 12:21]
  assign _T_422 = _T_420 | _T_421; // @[LZD.scala 49:16]
  assign _T_423 = ~ _T_421; // @[LZD.scala 49:27]
  assign _T_424 = _T_420 | _T_423; // @[LZD.scala 49:25]
  assign _T_425 = _T_412[0:0]; // @[LZD.scala 49:47]
  assign _T_426 = _T_419[0:0]; // @[LZD.scala 49:59]
  assign _T_427 = _T_420 ? _T_425 : _T_426; // @[LZD.scala 49:35]
  assign _T_429 = {_T_422,_T_424,_T_427}; // @[Cat.scala 29:58]
  assign _T_430 = _T_404[2]; // @[Shift.scala 12:21]
  assign _T_431 = _T_429[2]; // @[Shift.scala 12:21]
  assign _T_432 = _T_430 | _T_431; // @[LZD.scala 49:16]
  assign _T_433 = ~ _T_431; // @[LZD.scala 49:27]
  assign _T_434 = _T_430 | _T_433; // @[LZD.scala 49:25]
  assign _T_435 = _T_404[1:0]; // @[LZD.scala 49:47]
  assign _T_436 = _T_429[1:0]; // @[LZD.scala 49:59]
  assign _T_437 = _T_430 ? _T_435 : _T_436; // @[LZD.scala 49:35]
  assign _T_439 = {_T_432,_T_434,_T_437}; // @[Cat.scala 29:58]
  assign _T_440 = sumXor[7:0]; // @[LZD.scala 44:32]
  assign _T_441 = _T_440[7:4]; // @[LZD.scala 43:32]
  assign _T_442 = _T_441[3:2]; // @[LZD.scala 43:32]
  assign _T_443 = _T_442 != 2'h0; // @[LZD.scala 39:14]
  assign _T_444 = _T_442[1]; // @[LZD.scala 39:21]
  assign _T_445 = _T_442[0]; // @[LZD.scala 39:30]
  assign _T_446 = ~ _T_445; // @[LZD.scala 39:27]
  assign _T_447 = _T_444 | _T_446; // @[LZD.scala 39:25]
  assign _T_448 = {_T_443,_T_447}; // @[Cat.scala 29:58]
  assign _T_449 = _T_441[1:0]; // @[LZD.scala 44:32]
  assign _T_450 = _T_449 != 2'h0; // @[LZD.scala 39:14]
  assign _T_451 = _T_449[1]; // @[LZD.scala 39:21]
  assign _T_452 = _T_449[0]; // @[LZD.scala 39:30]
  assign _T_453 = ~ _T_452; // @[LZD.scala 39:27]
  assign _T_454 = _T_451 | _T_453; // @[LZD.scala 39:25]
  assign _T_455 = {_T_450,_T_454}; // @[Cat.scala 29:58]
  assign _T_456 = _T_448[1]; // @[Shift.scala 12:21]
  assign _T_457 = _T_455[1]; // @[Shift.scala 12:21]
  assign _T_458 = _T_456 | _T_457; // @[LZD.scala 49:16]
  assign _T_459 = ~ _T_457; // @[LZD.scala 49:27]
  assign _T_460 = _T_456 | _T_459; // @[LZD.scala 49:25]
  assign _T_461 = _T_448[0:0]; // @[LZD.scala 49:47]
  assign _T_462 = _T_455[0:0]; // @[LZD.scala 49:59]
  assign _T_463 = _T_456 ? _T_461 : _T_462; // @[LZD.scala 49:35]
  assign _T_465 = {_T_458,_T_460,_T_463}; // @[Cat.scala 29:58]
  assign _T_466 = _T_440[3:0]; // @[LZD.scala 44:32]
  assign _T_467 = _T_466[3:2]; // @[LZD.scala 43:32]
  assign _T_468 = _T_467 != 2'h0; // @[LZD.scala 39:14]
  assign _T_469 = _T_467[1]; // @[LZD.scala 39:21]
  assign _T_470 = _T_467[0]; // @[LZD.scala 39:30]
  assign _T_471 = ~ _T_470; // @[LZD.scala 39:27]
  assign _T_472 = _T_469 | _T_471; // @[LZD.scala 39:25]
  assign _T_473 = {_T_468,_T_472}; // @[Cat.scala 29:58]
  assign _T_474 = _T_466[1:0]; // @[LZD.scala 44:32]
  assign _T_475 = _T_474 != 2'h0; // @[LZD.scala 39:14]
  assign _T_476 = _T_474[1]; // @[LZD.scala 39:21]
  assign _T_477 = _T_474[0]; // @[LZD.scala 39:30]
  assign _T_478 = ~ _T_477; // @[LZD.scala 39:27]
  assign _T_479 = _T_476 | _T_478; // @[LZD.scala 39:25]
  assign _T_480 = {_T_475,_T_479}; // @[Cat.scala 29:58]
  assign _T_481 = _T_473[1]; // @[Shift.scala 12:21]
  assign _T_482 = _T_480[1]; // @[Shift.scala 12:21]
  assign _T_483 = _T_481 | _T_482; // @[LZD.scala 49:16]
  assign _T_484 = ~ _T_482; // @[LZD.scala 49:27]
  assign _T_485 = _T_481 | _T_484; // @[LZD.scala 49:25]
  assign _T_486 = _T_473[0:0]; // @[LZD.scala 49:47]
  assign _T_487 = _T_480[0:0]; // @[LZD.scala 49:59]
  assign _T_488 = _T_481 ? _T_486 : _T_487; // @[LZD.scala 49:35]
  assign _T_490 = {_T_483,_T_485,_T_488}; // @[Cat.scala 29:58]
  assign _T_491 = _T_465[2]; // @[Shift.scala 12:21]
  assign _T_492 = _T_490[2]; // @[Shift.scala 12:21]
  assign _T_493 = _T_491 | _T_492; // @[LZD.scala 49:16]
  assign _T_494 = ~ _T_492; // @[LZD.scala 49:27]
  assign _T_495 = _T_491 | _T_494; // @[LZD.scala 49:25]
  assign _T_496 = _T_465[1:0]; // @[LZD.scala 49:47]
  assign _T_497 = _T_490[1:0]; // @[LZD.scala 49:59]
  assign _T_498 = _T_491 ? _T_496 : _T_497; // @[LZD.scala 49:35]
  assign _T_500 = {_T_493,_T_495,_T_498}; // @[Cat.scala 29:58]
  assign _T_501 = _T_439[3]; // @[Shift.scala 12:21]
  assign _T_502 = _T_500[3]; // @[Shift.scala 12:21]
  assign _T_503 = _T_501 | _T_502; // @[LZD.scala 49:16]
  assign _T_504 = ~ _T_502; // @[LZD.scala 49:27]
  assign _T_505 = _T_501 | _T_504; // @[LZD.scala 49:25]
  assign _T_506 = _T_439[2:0]; // @[LZD.scala 49:47]
  assign _T_507 = _T_500[2:0]; // @[LZD.scala 49:59]
  assign _T_508 = _T_501 ? _T_506 : _T_507; // @[LZD.scala 49:35]
  assign sumLZD = {_T_503,_T_505,_T_508}; // @[Cat.scala 29:58]
  assign _T_510 = {1'h1,_T_503,_T_505,_T_508}; // @[Cat.scala 29:58]
  assign _T_511 = $signed(_T_510); // @[PositAdder.scala 41:38]
  assign _T_513 = $signed(_T_511) + $signed(6'sh2); // @[PositAdder.scala 41:45]
  assign scaleBias = $signed(_T_513); // @[PositAdder.scala 41:45]
  assign sumScale = $signed(greaterExp) + $signed(scaleBias); // @[PositAdder.scala 42:32]
  assign overflow = $signed(sumScale) > $signed(7'sh1a); // @[PositAdder.scala 43:30]
  assign normalShift = ~ sumLZD; // @[PositAdder.scala 44:22]
  assign _T_514 = signSumSig[14:0]; // @[PositAdder.scala 45:36]
  assign _T_515 = normalShift < 5'hf; // @[Shift.scala 16:24]
  assign _T_516 = normalShift[3:0]; // @[Shift.scala 17:37]
  assign _T_517 = _T_516[3]; // @[Shift.scala 12:21]
  assign _T_518 = _T_514[6:0]; // @[Shift.scala 64:52]
  assign _T_520 = {_T_518,8'h0}; // @[Cat.scala 29:58]
  assign _T_521 = _T_517 ? _T_520 : _T_514; // @[Shift.scala 64:27]
  assign _T_522 = _T_516[2:0]; // @[Shift.scala 66:70]
  assign _T_523 = _T_522[2]; // @[Shift.scala 12:21]
  assign _T_524 = _T_521[10:0]; // @[Shift.scala 64:52]
  assign _T_526 = {_T_524,4'h0}; // @[Cat.scala 29:58]
  assign _T_527 = _T_523 ? _T_526 : _T_521; // @[Shift.scala 64:27]
  assign _T_528 = _T_522[1:0]; // @[Shift.scala 66:70]
  assign _T_529 = _T_528[1]; // @[Shift.scala 12:21]
  assign _T_530 = _T_527[12:0]; // @[Shift.scala 64:52]
  assign _T_532 = {_T_530,2'h0}; // @[Cat.scala 29:58]
  assign _T_533 = _T_529 ? _T_532 : _T_527; // @[Shift.scala 64:27]
  assign _T_534 = _T_528[0:0]; // @[Shift.scala 66:70]
  assign _T_536 = _T_533[13:0]; // @[Shift.scala 64:52]
  assign _T_537 = {_T_536,1'h0}; // @[Cat.scala 29:58]
  assign _T_538 = _T_534 ? _T_537 : _T_533; // @[Shift.scala 64:27]
  assign shiftSig = _T_515 ? _T_538 : 15'h0; // @[Shift.scala 16:10]
  assign _T_539 = overflow ? $signed(7'sh1a) : $signed(sumScale); // @[PositAdder.scala 50:24]
  assign decS_fraction = shiftSig[14:4]; // @[PositAdder.scala 51:34]
  assign decS_isNaR = decA_isNaR | decB_isNaR; // @[PositAdder.scala 52:32]
  assign _T_542 = signSumSig != 17'h0; // @[PositAdder.scala 53:33]
  assign _T_543 = ~ _T_542; // @[PositAdder.scala 53:21]
  assign _T_544 = decA_isZero & decB_isZero; // @[PositAdder.scala 53:52]
  assign decS_isZero = _T_543 | _T_544; // @[PositAdder.scala 53:37]
  assign _T_546 = shiftSig[3:2]; // @[PositAdder.scala 54:33]
  assign _T_547 = shiftSig[1]; // @[PositAdder.scala 54:49]
  assign _T_548 = shiftSig[0]; // @[PositAdder.scala 54:63]
  assign _T_549 = _T_547 | _T_548; // @[PositAdder.scala 54:53]
  assign _GEN_4 = _T_539[5:0]; // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  assign decS_scale = $signed(_GEN_4); // @[PositAdder.scala 47:25 PositAdder.scala 50:18]
  assign _T_552 = decS_scale[0]; // @[convert.scala 46:61]
  assign _T_553 = ~ _T_552; // @[convert.scala 46:52]
  assign _T_555 = sumSign ? _T_553 : _T_552; // @[convert.scala 46:42]
  assign _T_556 = decS_scale[5:1]; // @[convert.scala 48:34]
  assign _T_557 = _T_556[4:4]; // @[convert.scala 49:36]
  assign _T_559 = ~ _T_556; // @[convert.scala 50:36]
  assign _T_560 = $signed(_T_559); // @[convert.scala 50:36]
  assign _T_561 = _T_557 ? $signed(_T_560) : $signed(_T_556); // @[convert.scala 50:28]
  assign _T_562 = _T_557 ^ sumSign; // @[convert.scala 51:31]
  assign _T_563 = ~ _T_562; // @[convert.scala 52:43]
  assign _T_567 = {_T_563,_T_562,_T_555,decS_fraction,_T_546,_T_549}; // @[Cat.scala 29:58]
  assign _T_568 = $unsigned(_T_561); // @[Shift.scala 39:17]
  assign _T_569 = _T_568 < 5'h11; // @[Shift.scala 39:24]
  assign _T_571 = _T_567[16:16]; // @[Shift.scala 90:30]
  assign _T_572 = _T_567[15:0]; // @[Shift.scala 90:48]
  assign _T_573 = _T_572 != 16'h0; // @[Shift.scala 90:57]
  assign _T_574 = _T_571 | _T_573; // @[Shift.scala 90:39]
  assign _T_575 = _T_568[4]; // @[Shift.scala 12:21]
  assign _T_576 = _T_567[16]; // @[Shift.scala 12:21]
  assign _T_578 = _T_576 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_579 = {_T_578,_T_574}; // @[Cat.scala 29:58]
  assign _T_580 = _T_575 ? _T_579 : _T_567; // @[Shift.scala 91:22]
  assign _T_581 = _T_568[3:0]; // @[Shift.scala 92:77]
  assign _T_582 = _T_580[16:8]; // @[Shift.scala 90:30]
  assign _T_583 = _T_580[7:0]; // @[Shift.scala 90:48]
  assign _T_584 = _T_583 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{8'd0}, _T_584}; // @[Shift.scala 90:39]
  assign _T_585 = _T_582 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_586 = _T_581[3]; // @[Shift.scala 12:21]
  assign _T_587 = _T_580[16]; // @[Shift.scala 12:21]
  assign _T_589 = _T_587 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_590 = {_T_589,_T_585}; // @[Cat.scala 29:58]
  assign _T_591 = _T_586 ? _T_590 : _T_580; // @[Shift.scala 91:22]
  assign _T_592 = _T_581[2:0]; // @[Shift.scala 92:77]
  assign _T_593 = _T_591[16:4]; // @[Shift.scala 90:30]
  assign _T_594 = _T_591[3:0]; // @[Shift.scala 90:48]
  assign _T_595 = _T_594 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{12'd0}, _T_595}; // @[Shift.scala 90:39]
  assign _T_596 = _T_593 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_597 = _T_592[2]; // @[Shift.scala 12:21]
  assign _T_598 = _T_591[16]; // @[Shift.scala 12:21]
  assign _T_600 = _T_598 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_601 = {_T_600,_T_596}; // @[Cat.scala 29:58]
  assign _T_602 = _T_597 ? _T_601 : _T_591; // @[Shift.scala 91:22]
  assign _T_603 = _T_592[1:0]; // @[Shift.scala 92:77]
  assign _T_604 = _T_602[16:2]; // @[Shift.scala 90:30]
  assign _T_605 = _T_602[1:0]; // @[Shift.scala 90:48]
  assign _T_606 = _T_605 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{14'd0}, _T_606}; // @[Shift.scala 90:39]
  assign _T_607 = _T_604 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_608 = _T_603[1]; // @[Shift.scala 12:21]
  assign _T_609 = _T_602[16]; // @[Shift.scala 12:21]
  assign _T_611 = _T_609 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_612 = {_T_611,_T_607}; // @[Cat.scala 29:58]
  assign _T_613 = _T_608 ? _T_612 : _T_602; // @[Shift.scala 91:22]
  assign _T_614 = _T_603[0:0]; // @[Shift.scala 92:77]
  assign _T_615 = _T_613[16:1]; // @[Shift.scala 90:30]
  assign _T_616 = _T_613[0:0]; // @[Shift.scala 90:48]
  assign _GEN_8 = {{15'd0}, _T_616}; // @[Shift.scala 90:39]
  assign _T_618 = _T_615 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_620 = _T_613[16]; // @[Shift.scala 12:21]
  assign _T_621 = {_T_620,_T_618}; // @[Cat.scala 29:58]
  assign _T_622 = _T_614 ? _T_621 : _T_613; // @[Shift.scala 91:22]
  assign _T_625 = _T_576 ? 17'h1ffff : 17'h0; // @[Bitwise.scala 71:12]
  assign _T_626 = _T_569 ? _T_622 : _T_625; // @[Shift.scala 39:10]
  assign _T_627 = _T_626[3]; // @[convert.scala 55:31]
  assign _T_628 = _T_626[2]; // @[convert.scala 56:31]
  assign _T_629 = _T_626[1]; // @[convert.scala 57:31]
  assign _T_630 = _T_626[0]; // @[convert.scala 58:31]
  assign _T_631 = _T_626[16:3]; // @[convert.scala 59:69]
  assign _T_632 = _T_631 != 14'h0; // @[convert.scala 59:81]
  assign _T_633 = ~ _T_632; // @[convert.scala 59:50]
  assign _T_635 = _T_631 == 14'h3fff; // @[convert.scala 60:81]
  assign _T_636 = _T_627 | _T_629; // @[convert.scala 61:44]
  assign _T_637 = _T_636 | _T_630; // @[convert.scala 61:52]
  assign _T_638 = _T_628 & _T_637; // @[convert.scala 61:36]
  assign _T_639 = ~ _T_635; // @[convert.scala 62:63]
  assign _T_640 = _T_639 & _T_638; // @[convert.scala 62:103]
  assign _T_641 = _T_633 | _T_640; // @[convert.scala 62:60]
  assign _GEN_9 = {{13'd0}, _T_641}; // @[convert.scala 63:56]
  assign _T_644 = _T_631 + _GEN_9; // @[convert.scala 63:56]
  assign _T_645 = {sumSign,_T_644}; // @[Cat.scala 29:58]
  assign _T_647 = decS_isZero ? 15'h0 : _T_645; // @[Mux.scala 87:16]
  assign io_S = decS_isNaR ? 15'h4000 : _T_647; // @[PositAdder.scala 56:8]
endmodule
