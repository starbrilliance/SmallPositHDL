module PositFMA13_1(
  input         clock,
  input         reset,
  input         io_inValid,
  input  [1:0]  io_fmaOp,
  input  [12:0] io_A,
  input  [12:0] io_B,
  input  [12:0] io_C,
  output [12:0] io_F,
  output        io_outValid
);
  wire  _T; // @[PositFMA.scala 47:36]
  wire [12:0] _T_2; // @[Bitwise.scala 71:12]
  wire [12:0] _T_3; // @[PositFMA.scala 47:41]
  wire [12:0] _GEN_10; // @[PositFMA.scala 47:49]
  wire [12:0] realA; // @[PositFMA.scala 47:49]
  wire  _T_6; // @[PositFMA.scala 48:36]
  wire [12:0] _T_8; // @[Bitwise.scala 71:12]
  wire [12:0] _T_9; // @[PositFMA.scala 48:41]
  wire [12:0] _GEN_11; // @[PositFMA.scala 48:49]
  wire [12:0] realC; // @[PositFMA.scala 48:49]
  wire  _T_13; // @[convert.scala 18:24]
  wire  _T_14; // @[convert.scala 18:40]
  wire  _T_15; // @[convert.scala 18:36]
  wire [10:0] _T_16; // @[convert.scala 19:24]
  wire [10:0] _T_17; // @[convert.scala 19:43]
  wire [10:0] _T_18; // @[convert.scala 19:39]
  wire [7:0] _T_19; // @[LZD.scala 43:32]
  wire [3:0] _T_20; // @[LZD.scala 43:32]
  wire [1:0] _T_21; // @[LZD.scala 43:32]
  wire  _T_22; // @[LZD.scala 39:14]
  wire  _T_23; // @[LZD.scala 39:21]
  wire  _T_24; // @[LZD.scala 39:30]
  wire  _T_25; // @[LZD.scala 39:27]
  wire  _T_26; // @[LZD.scala 39:25]
  wire [1:0] _T_27; // @[Cat.scala 29:58]
  wire [1:0] _T_28; // @[LZD.scala 44:32]
  wire  _T_29; // @[LZD.scala 39:14]
  wire  _T_30; // @[LZD.scala 39:21]
  wire  _T_31; // @[LZD.scala 39:30]
  wire  _T_32; // @[LZD.scala 39:27]
  wire  _T_33; // @[LZD.scala 39:25]
  wire [1:0] _T_34; // @[Cat.scala 29:58]
  wire  _T_35; // @[Shift.scala 12:21]
  wire  _T_36; // @[Shift.scala 12:21]
  wire  _T_37; // @[LZD.scala 49:16]
  wire  _T_38; // @[LZD.scala 49:27]
  wire  _T_39; // @[LZD.scala 49:25]
  wire  _T_40; // @[LZD.scala 49:47]
  wire  _T_41; // @[LZD.scala 49:59]
  wire  _T_42; // @[LZD.scala 49:35]
  wire [2:0] _T_44; // @[Cat.scala 29:58]
  wire [3:0] _T_45; // @[LZD.scala 44:32]
  wire [1:0] _T_46; // @[LZD.scala 43:32]
  wire  _T_47; // @[LZD.scala 39:14]
  wire  _T_48; // @[LZD.scala 39:21]
  wire  _T_49; // @[LZD.scala 39:30]
  wire  _T_50; // @[LZD.scala 39:27]
  wire  _T_51; // @[LZD.scala 39:25]
  wire [1:0] _T_52; // @[Cat.scala 29:58]
  wire [1:0] _T_53; // @[LZD.scala 44:32]
  wire  _T_54; // @[LZD.scala 39:14]
  wire  _T_55; // @[LZD.scala 39:21]
  wire  _T_56; // @[LZD.scala 39:30]
  wire  _T_57; // @[LZD.scala 39:27]
  wire  _T_58; // @[LZD.scala 39:25]
  wire [1:0] _T_59; // @[Cat.scala 29:58]
  wire  _T_60; // @[Shift.scala 12:21]
  wire  _T_61; // @[Shift.scala 12:21]
  wire  _T_62; // @[LZD.scala 49:16]
  wire  _T_63; // @[LZD.scala 49:27]
  wire  _T_64; // @[LZD.scala 49:25]
  wire  _T_65; // @[LZD.scala 49:47]
  wire  _T_66; // @[LZD.scala 49:59]
  wire  _T_67; // @[LZD.scala 49:35]
  wire [2:0] _T_69; // @[Cat.scala 29:58]
  wire  _T_70; // @[Shift.scala 12:21]
  wire  _T_71; // @[Shift.scala 12:21]
  wire  _T_72; // @[LZD.scala 49:16]
  wire  _T_73; // @[LZD.scala 49:27]
  wire  _T_74; // @[LZD.scala 49:25]
  wire [1:0] _T_75; // @[LZD.scala 49:47]
  wire [1:0] _T_76; // @[LZD.scala 49:59]
  wire [1:0] _T_77; // @[LZD.scala 49:35]
  wire [3:0] _T_79; // @[Cat.scala 29:58]
  wire [2:0] _T_80; // @[LZD.scala 44:32]
  wire [1:0] _T_81; // @[LZD.scala 43:32]
  wire  _T_82; // @[LZD.scala 39:14]
  wire  _T_83; // @[LZD.scala 39:21]
  wire  _T_84; // @[LZD.scala 39:30]
  wire  _T_85; // @[LZD.scala 39:27]
  wire  _T_86; // @[LZD.scala 39:25]
  wire [1:0] _T_87; // @[Cat.scala 29:58]
  wire  _T_88; // @[LZD.scala 44:32]
  wire  _T_90; // @[Shift.scala 12:21]
  wire  _T_92; // @[LZD.scala 55:32]
  wire  _T_93; // @[LZD.scala 55:20]
  wire  _T_95; // @[Shift.scala 12:21]
  wire [2:0] _T_97; // @[Cat.scala 29:58]
  wire [2:0] _T_98; // @[LZD.scala 55:32]
  wire [2:0] _T_99; // @[LZD.scala 55:20]
  wire [3:0] _T_100; // @[Cat.scala 29:58]
  wire [3:0] _T_101; // @[convert.scala 21:22]
  wire [9:0] _T_102; // @[convert.scala 22:36]
  wire  _T_103; // @[Shift.scala 16:24]
  wire  _T_105; // @[Shift.scala 12:21]
  wire [1:0] _T_106; // @[Shift.scala 64:52]
  wire [9:0] _T_108; // @[Cat.scala 29:58]
  wire [9:0] _T_109; // @[Shift.scala 64:27]
  wire [2:0] _T_110; // @[Shift.scala 66:70]
  wire  _T_111; // @[Shift.scala 12:21]
  wire [5:0] _T_112; // @[Shift.scala 64:52]
  wire [9:0] _T_114; // @[Cat.scala 29:58]
  wire [9:0] _T_115; // @[Shift.scala 64:27]
  wire [1:0] _T_116; // @[Shift.scala 66:70]
  wire  _T_117; // @[Shift.scala 12:21]
  wire [7:0] _T_118; // @[Shift.scala 64:52]
  wire [9:0] _T_120; // @[Cat.scala 29:58]
  wire [9:0] _T_121; // @[Shift.scala 64:27]
  wire  _T_122; // @[Shift.scala 66:70]
  wire [8:0] _T_124; // @[Shift.scala 64:52]
  wire [9:0] _T_125; // @[Cat.scala 29:58]
  wire [9:0] _T_126; // @[Shift.scala 64:27]
  wire [9:0] _T_127; // @[Shift.scala 16:10]
  wire  _T_128; // @[convert.scala 23:34]
  wire [8:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_130; // @[convert.scala 25:26]
  wire [3:0] _T_132; // @[convert.scala 25:42]
  wire  _T_135; // @[convert.scala 26:67]
  wire  _T_136; // @[convert.scala 26:51]
  wire [5:0] _T_137; // @[Cat.scala 29:58]
  wire [11:0] _T_139; // @[convert.scala 29:56]
  wire  _T_140; // @[convert.scala 29:60]
  wire  _T_141; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_144; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_153; // @[convert.scala 18:24]
  wire  _T_154; // @[convert.scala 18:40]
  wire  _T_155; // @[convert.scala 18:36]
  wire [10:0] _T_156; // @[convert.scala 19:24]
  wire [10:0] _T_157; // @[convert.scala 19:43]
  wire [10:0] _T_158; // @[convert.scala 19:39]
  wire [7:0] _T_159; // @[LZD.scala 43:32]
  wire [3:0] _T_160; // @[LZD.scala 43:32]
  wire [1:0] _T_161; // @[LZD.scala 43:32]
  wire  _T_162; // @[LZD.scala 39:14]
  wire  _T_163; // @[LZD.scala 39:21]
  wire  _T_164; // @[LZD.scala 39:30]
  wire  _T_165; // @[LZD.scala 39:27]
  wire  _T_166; // @[LZD.scala 39:25]
  wire [1:0] _T_167; // @[Cat.scala 29:58]
  wire [1:0] _T_168; // @[LZD.scala 44:32]
  wire  _T_169; // @[LZD.scala 39:14]
  wire  _T_170; // @[LZD.scala 39:21]
  wire  _T_171; // @[LZD.scala 39:30]
  wire  _T_172; // @[LZD.scala 39:27]
  wire  _T_173; // @[LZD.scala 39:25]
  wire [1:0] _T_174; // @[Cat.scala 29:58]
  wire  _T_175; // @[Shift.scala 12:21]
  wire  _T_176; // @[Shift.scala 12:21]
  wire  _T_177; // @[LZD.scala 49:16]
  wire  _T_178; // @[LZD.scala 49:27]
  wire  _T_179; // @[LZD.scala 49:25]
  wire  _T_180; // @[LZD.scala 49:47]
  wire  _T_181; // @[LZD.scala 49:59]
  wire  _T_182; // @[LZD.scala 49:35]
  wire [2:0] _T_184; // @[Cat.scala 29:58]
  wire [3:0] _T_185; // @[LZD.scala 44:32]
  wire [1:0] _T_186; // @[LZD.scala 43:32]
  wire  _T_187; // @[LZD.scala 39:14]
  wire  _T_188; // @[LZD.scala 39:21]
  wire  _T_189; // @[LZD.scala 39:30]
  wire  _T_190; // @[LZD.scala 39:27]
  wire  _T_191; // @[LZD.scala 39:25]
  wire [1:0] _T_192; // @[Cat.scala 29:58]
  wire [1:0] _T_193; // @[LZD.scala 44:32]
  wire  _T_194; // @[LZD.scala 39:14]
  wire  _T_195; // @[LZD.scala 39:21]
  wire  _T_196; // @[LZD.scala 39:30]
  wire  _T_197; // @[LZD.scala 39:27]
  wire  _T_198; // @[LZD.scala 39:25]
  wire [1:0] _T_199; // @[Cat.scala 29:58]
  wire  _T_200; // @[Shift.scala 12:21]
  wire  _T_201; // @[Shift.scala 12:21]
  wire  _T_202; // @[LZD.scala 49:16]
  wire  _T_203; // @[LZD.scala 49:27]
  wire  _T_204; // @[LZD.scala 49:25]
  wire  _T_205; // @[LZD.scala 49:47]
  wire  _T_206; // @[LZD.scala 49:59]
  wire  _T_207; // @[LZD.scala 49:35]
  wire [2:0] _T_209; // @[Cat.scala 29:58]
  wire  _T_210; // @[Shift.scala 12:21]
  wire  _T_211; // @[Shift.scala 12:21]
  wire  _T_212; // @[LZD.scala 49:16]
  wire  _T_213; // @[LZD.scala 49:27]
  wire  _T_214; // @[LZD.scala 49:25]
  wire [1:0] _T_215; // @[LZD.scala 49:47]
  wire [1:0] _T_216; // @[LZD.scala 49:59]
  wire [1:0] _T_217; // @[LZD.scala 49:35]
  wire [3:0] _T_219; // @[Cat.scala 29:58]
  wire [2:0] _T_220; // @[LZD.scala 44:32]
  wire [1:0] _T_221; // @[LZD.scala 43:32]
  wire  _T_222; // @[LZD.scala 39:14]
  wire  _T_223; // @[LZD.scala 39:21]
  wire  _T_224; // @[LZD.scala 39:30]
  wire  _T_225; // @[LZD.scala 39:27]
  wire  _T_226; // @[LZD.scala 39:25]
  wire [1:0] _T_227; // @[Cat.scala 29:58]
  wire  _T_228; // @[LZD.scala 44:32]
  wire  _T_230; // @[Shift.scala 12:21]
  wire  _T_232; // @[LZD.scala 55:32]
  wire  _T_233; // @[LZD.scala 55:20]
  wire  _T_235; // @[Shift.scala 12:21]
  wire [2:0] _T_237; // @[Cat.scala 29:58]
  wire [2:0] _T_238; // @[LZD.scala 55:32]
  wire [2:0] _T_239; // @[LZD.scala 55:20]
  wire [3:0] _T_240; // @[Cat.scala 29:58]
  wire [3:0] _T_241; // @[convert.scala 21:22]
  wire [9:0] _T_242; // @[convert.scala 22:36]
  wire  _T_243; // @[Shift.scala 16:24]
  wire  _T_245; // @[Shift.scala 12:21]
  wire [1:0] _T_246; // @[Shift.scala 64:52]
  wire [9:0] _T_248; // @[Cat.scala 29:58]
  wire [9:0] _T_249; // @[Shift.scala 64:27]
  wire [2:0] _T_250; // @[Shift.scala 66:70]
  wire  _T_251; // @[Shift.scala 12:21]
  wire [5:0] _T_252; // @[Shift.scala 64:52]
  wire [9:0] _T_254; // @[Cat.scala 29:58]
  wire [9:0] _T_255; // @[Shift.scala 64:27]
  wire [1:0] _T_256; // @[Shift.scala 66:70]
  wire  _T_257; // @[Shift.scala 12:21]
  wire [7:0] _T_258; // @[Shift.scala 64:52]
  wire [9:0] _T_260; // @[Cat.scala 29:58]
  wire [9:0] _T_261; // @[Shift.scala 64:27]
  wire  _T_262; // @[Shift.scala 66:70]
  wire [8:0] _T_264; // @[Shift.scala 64:52]
  wire [9:0] _T_265; // @[Cat.scala 29:58]
  wire [9:0] _T_266; // @[Shift.scala 64:27]
  wire [9:0] _T_267; // @[Shift.scala 16:10]
  wire  _T_268; // @[convert.scala 23:34]
  wire [8:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_270; // @[convert.scala 25:26]
  wire [3:0] _T_272; // @[convert.scala 25:42]
  wire  _T_275; // @[convert.scala 26:67]
  wire  _T_276; // @[convert.scala 26:51]
  wire [5:0] _T_277; // @[Cat.scala 29:58]
  wire [11:0] _T_279; // @[convert.scala 29:56]
  wire  _T_280; // @[convert.scala 29:60]
  wire  _T_281; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_284; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_293; // @[convert.scala 18:24]
  wire  _T_294; // @[convert.scala 18:40]
  wire  _T_295; // @[convert.scala 18:36]
  wire [10:0] _T_296; // @[convert.scala 19:24]
  wire [10:0] _T_297; // @[convert.scala 19:43]
  wire [10:0] _T_298; // @[convert.scala 19:39]
  wire [7:0] _T_299; // @[LZD.scala 43:32]
  wire [3:0] _T_300; // @[LZD.scala 43:32]
  wire [1:0] _T_301; // @[LZD.scala 43:32]
  wire  _T_302; // @[LZD.scala 39:14]
  wire  _T_303; // @[LZD.scala 39:21]
  wire  _T_304; // @[LZD.scala 39:30]
  wire  _T_305; // @[LZD.scala 39:27]
  wire  _T_306; // @[LZD.scala 39:25]
  wire [1:0] _T_307; // @[Cat.scala 29:58]
  wire [1:0] _T_308; // @[LZD.scala 44:32]
  wire  _T_309; // @[LZD.scala 39:14]
  wire  _T_310; // @[LZD.scala 39:21]
  wire  _T_311; // @[LZD.scala 39:30]
  wire  _T_312; // @[LZD.scala 39:27]
  wire  _T_313; // @[LZD.scala 39:25]
  wire [1:0] _T_314; // @[Cat.scala 29:58]
  wire  _T_315; // @[Shift.scala 12:21]
  wire  _T_316; // @[Shift.scala 12:21]
  wire  _T_317; // @[LZD.scala 49:16]
  wire  _T_318; // @[LZD.scala 49:27]
  wire  _T_319; // @[LZD.scala 49:25]
  wire  _T_320; // @[LZD.scala 49:47]
  wire  _T_321; // @[LZD.scala 49:59]
  wire  _T_322; // @[LZD.scala 49:35]
  wire [2:0] _T_324; // @[Cat.scala 29:58]
  wire [3:0] _T_325; // @[LZD.scala 44:32]
  wire [1:0] _T_326; // @[LZD.scala 43:32]
  wire  _T_327; // @[LZD.scala 39:14]
  wire  _T_328; // @[LZD.scala 39:21]
  wire  _T_329; // @[LZD.scala 39:30]
  wire  _T_330; // @[LZD.scala 39:27]
  wire  _T_331; // @[LZD.scala 39:25]
  wire [1:0] _T_332; // @[Cat.scala 29:58]
  wire [1:0] _T_333; // @[LZD.scala 44:32]
  wire  _T_334; // @[LZD.scala 39:14]
  wire  _T_335; // @[LZD.scala 39:21]
  wire  _T_336; // @[LZD.scala 39:30]
  wire  _T_337; // @[LZD.scala 39:27]
  wire  _T_338; // @[LZD.scala 39:25]
  wire [1:0] _T_339; // @[Cat.scala 29:58]
  wire  _T_340; // @[Shift.scala 12:21]
  wire  _T_341; // @[Shift.scala 12:21]
  wire  _T_342; // @[LZD.scala 49:16]
  wire  _T_343; // @[LZD.scala 49:27]
  wire  _T_344; // @[LZD.scala 49:25]
  wire  _T_345; // @[LZD.scala 49:47]
  wire  _T_346; // @[LZD.scala 49:59]
  wire  _T_347; // @[LZD.scala 49:35]
  wire [2:0] _T_349; // @[Cat.scala 29:58]
  wire  _T_350; // @[Shift.scala 12:21]
  wire  _T_351; // @[Shift.scala 12:21]
  wire  _T_352; // @[LZD.scala 49:16]
  wire  _T_353; // @[LZD.scala 49:27]
  wire  _T_354; // @[LZD.scala 49:25]
  wire [1:0] _T_355; // @[LZD.scala 49:47]
  wire [1:0] _T_356; // @[LZD.scala 49:59]
  wire [1:0] _T_357; // @[LZD.scala 49:35]
  wire [3:0] _T_359; // @[Cat.scala 29:58]
  wire [2:0] _T_360; // @[LZD.scala 44:32]
  wire [1:0] _T_361; // @[LZD.scala 43:32]
  wire  _T_362; // @[LZD.scala 39:14]
  wire  _T_363; // @[LZD.scala 39:21]
  wire  _T_364; // @[LZD.scala 39:30]
  wire  _T_365; // @[LZD.scala 39:27]
  wire  _T_366; // @[LZD.scala 39:25]
  wire [1:0] _T_367; // @[Cat.scala 29:58]
  wire  _T_368; // @[LZD.scala 44:32]
  wire  _T_370; // @[Shift.scala 12:21]
  wire  _T_372; // @[LZD.scala 55:32]
  wire  _T_373; // @[LZD.scala 55:20]
  wire  _T_375; // @[Shift.scala 12:21]
  wire [2:0] _T_377; // @[Cat.scala 29:58]
  wire [2:0] _T_378; // @[LZD.scala 55:32]
  wire [2:0] _T_379; // @[LZD.scala 55:20]
  wire [3:0] _T_380; // @[Cat.scala 29:58]
  wire [3:0] _T_381; // @[convert.scala 21:22]
  wire [9:0] _T_382; // @[convert.scala 22:36]
  wire  _T_383; // @[Shift.scala 16:24]
  wire  _T_385; // @[Shift.scala 12:21]
  wire [1:0] _T_386; // @[Shift.scala 64:52]
  wire [9:0] _T_388; // @[Cat.scala 29:58]
  wire [9:0] _T_389; // @[Shift.scala 64:27]
  wire [2:0] _T_390; // @[Shift.scala 66:70]
  wire  _T_391; // @[Shift.scala 12:21]
  wire [5:0] _T_392; // @[Shift.scala 64:52]
  wire [9:0] _T_394; // @[Cat.scala 29:58]
  wire [9:0] _T_395; // @[Shift.scala 64:27]
  wire [1:0] _T_396; // @[Shift.scala 66:70]
  wire  _T_397; // @[Shift.scala 12:21]
  wire [7:0] _T_398; // @[Shift.scala 64:52]
  wire [9:0] _T_400; // @[Cat.scala 29:58]
  wire [9:0] _T_401; // @[Shift.scala 64:27]
  wire  _T_402; // @[Shift.scala 66:70]
  wire [8:0] _T_404; // @[Shift.scala 64:52]
  wire [9:0] _T_405; // @[Cat.scala 29:58]
  wire [9:0] _T_406; // @[Shift.scala 64:27]
  wire [9:0] _T_407; // @[Shift.scala 16:10]
  wire  _T_408; // @[convert.scala 23:34]
  wire [8:0] decC_fraction; // @[convert.scala 24:34]
  wire  _T_410; // @[convert.scala 25:26]
  wire [3:0] _T_412; // @[convert.scala 25:42]
  wire  _T_415; // @[convert.scala 26:67]
  wire  _T_416; // @[convert.scala 26:51]
  wire [5:0] _T_417; // @[Cat.scala 29:58]
  wire [11:0] _T_419; // @[convert.scala 29:56]
  wire  _T_420; // @[convert.scala 29:60]
  wire  _T_421; // @[convert.scala 29:41]
  wire  decC_isNaR; // @[convert.scala 29:39]
  wire  _T_424; // @[convert.scala 30:19]
  wire  decC_isZero; // @[convert.scala 30:41]
  wire [5:0] decC_scale; // @[convert.scala 32:24]
  wire  _T_432; // @[PositFMA.scala 58:30]
  wire  outIsNaR; // @[PositFMA.scala 58:44]
  wire  _T_433; // @[PositFMA.scala 59:34]
  wire  _T_434; // @[PositFMA.scala 59:47]
  wire  _T_435; // @[PositFMA.scala 59:45]
  wire [10:0] _T_437; // @[Cat.scala 29:58]
  wire [10:0] sigA; // @[PositFMA.scala 59:76]
  wire  _T_438; // @[PositFMA.scala 60:34]
  wire  _T_439; // @[PositFMA.scala 60:47]
  wire  _T_440; // @[PositFMA.scala 60:45]
  wire [10:0] _T_442; // @[Cat.scala 29:58]
  wire [10:0] sigB; // @[PositFMA.scala 60:76]
  wire [21:0] _T_443; // @[PositFMA.scala 61:25]
  wire [21:0] sigP; // @[PositFMA.scala 61:33]
  wire [18:0] _T_444; // @[PositFMA.scala 62:29]
  wire  _T_445; // @[PositFMA.scala 62:33]
  wire  eqTwo; // @[PositFMA.scala 62:19]
  wire  _T_446; // @[PositFMA.scala 64:29]
  wire  _T_447; // @[PositFMA.scala 64:56]
  wire  _T_448; // @[PositFMA.scala 64:51]
  wire  _T_449; // @[PositFMA.scala 64:49]
  wire  eqFour; // @[PositFMA.scala 64:76]
  wire  _T_450; // @[PositFMA.scala 66:23]
  wire  geTwo; // @[PositFMA.scala 66:43]
  wire [1:0] _T_452; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositFMA.scala 67:38]
  wire  mulSign; // @[PositFMA.scala 68:28]
  wire [6:0] _T_453; // @[PositFMA.scala 70:30]
  wire [6:0] _GEN_12; // @[PositFMA.scala 70:44]
  wire [6:0] _T_455; // @[PositFMA.scala 70:44]
  wire [6:0] mulScale; // @[PositFMA.scala 70:44]
  wire [19:0] _T_456; // @[PositFMA.scala 73:29]
  wire [18:0] _T_457; // @[PositFMA.scala 74:29]
  wire [19:0] _T_458; // @[PositFMA.scala 74:48]
  wire [19:0] mulSigTmp; // @[PositFMA.scala 71:22]
  wire  _T_460; // @[PositFMA.scala 78:39]
  wire  _T_461; // @[PositFMA.scala 78:43]
  wire [18:0] _T_462; // @[PositFMA.scala 79:39]
  wire [20:0] mulSig; // @[Cat.scala 29:58]
  reg  outIsNaR_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg [20:0] mulSig_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [8:0] addFrac_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [6:0] mulScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [5:0] addScale_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  addSign_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  addZero_phase2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  inValid_phase2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_7;
  wire  _T_488; // @[PositFMA.scala 108:29]
  wire  _T_489; // @[PositFMA.scala 108:47]
  wire  _T_490; // @[PositFMA.scala 108:45]
  wire [20:0] extAddSig; // @[Cat.scala 29:58]
  wire [6:0] _GEN_13; // @[PositFMA.scala 112:39]
  wire  mulGreater; // @[PositFMA.scala 112:39]
  wire [6:0] greaterScale; // @[PositFMA.scala 113:26]
  wire [6:0] smallerScale; // @[PositFMA.scala 114:26]
  wire [6:0] _T_494; // @[PositFMA.scala 115:36]
  wire [6:0] scaleDiff; // @[PositFMA.scala 115:36]
  wire [20:0] greaterSig; // @[PositFMA.scala 116:26]
  wire [20:0] smallerSigTmp; // @[PositFMA.scala 117:26]
  wire [6:0] _T_495; // @[PositFMA.scala 118:69]
  wire  _T_496; // @[Shift.scala 39:24]
  wire [4:0] _T_497; // @[Shift.scala 40:44]
  wire [4:0] _T_498; // @[Shift.scala 90:30]
  wire [15:0] _T_499; // @[Shift.scala 90:48]
  wire  _T_500; // @[Shift.scala 90:57]
  wire [4:0] _GEN_14; // @[Shift.scala 90:39]
  wire [4:0] _T_501; // @[Shift.scala 90:39]
  wire  _T_502; // @[Shift.scala 12:21]
  wire  _T_503; // @[Shift.scala 12:21]
  wire [15:0] _T_505; // @[Bitwise.scala 71:12]
  wire [20:0] _T_506; // @[Cat.scala 29:58]
  wire [20:0] _T_507; // @[Shift.scala 91:22]
  wire [3:0] _T_508; // @[Shift.scala 92:77]
  wire [12:0] _T_509; // @[Shift.scala 90:30]
  wire [7:0] _T_510; // @[Shift.scala 90:48]
  wire  _T_511; // @[Shift.scala 90:57]
  wire [12:0] _GEN_15; // @[Shift.scala 90:39]
  wire [12:0] _T_512; // @[Shift.scala 90:39]
  wire  _T_513; // @[Shift.scala 12:21]
  wire  _T_514; // @[Shift.scala 12:21]
  wire [7:0] _T_516; // @[Bitwise.scala 71:12]
  wire [20:0] _T_517; // @[Cat.scala 29:58]
  wire [20:0] _T_518; // @[Shift.scala 91:22]
  wire [2:0] _T_519; // @[Shift.scala 92:77]
  wire [16:0] _T_520; // @[Shift.scala 90:30]
  wire [3:0] _T_521; // @[Shift.scala 90:48]
  wire  _T_522; // @[Shift.scala 90:57]
  wire [16:0] _GEN_16; // @[Shift.scala 90:39]
  wire [16:0] _T_523; // @[Shift.scala 90:39]
  wire  _T_524; // @[Shift.scala 12:21]
  wire  _T_525; // @[Shift.scala 12:21]
  wire [3:0] _T_527; // @[Bitwise.scala 71:12]
  wire [20:0] _T_528; // @[Cat.scala 29:58]
  wire [20:0] _T_529; // @[Shift.scala 91:22]
  wire [1:0] _T_530; // @[Shift.scala 92:77]
  wire [18:0] _T_531; // @[Shift.scala 90:30]
  wire [1:0] _T_532; // @[Shift.scala 90:48]
  wire  _T_533; // @[Shift.scala 90:57]
  wire [18:0] _GEN_17; // @[Shift.scala 90:39]
  wire [18:0] _T_534; // @[Shift.scala 90:39]
  wire  _T_535; // @[Shift.scala 12:21]
  wire  _T_536; // @[Shift.scala 12:21]
  wire [1:0] _T_538; // @[Bitwise.scala 71:12]
  wire [20:0] _T_539; // @[Cat.scala 29:58]
  wire [20:0] _T_540; // @[Shift.scala 91:22]
  wire  _T_541; // @[Shift.scala 92:77]
  wire [19:0] _T_542; // @[Shift.scala 90:30]
  wire  _T_543; // @[Shift.scala 90:48]
  wire [19:0] _GEN_18; // @[Shift.scala 90:39]
  wire [19:0] _T_545; // @[Shift.scala 90:39]
  wire  _T_547; // @[Shift.scala 12:21]
  wire [20:0] _T_548; // @[Cat.scala 29:58]
  wire [20:0] _T_549; // @[Shift.scala 91:22]
  wire [20:0] _T_552; // @[Bitwise.scala 71:12]
  wire [20:0] smallerSig; // @[Shift.scala 39:10]
  wire [21:0] rawSumSig; // @[PositFMA.scala 119:34]
  wire  _T_553; // @[PositFMA.scala 120:42]
  wire  _T_554; // @[PositFMA.scala 120:46]
  wire  _T_555; // @[PositFMA.scala 120:79]
  wire  sumSign; // @[PositFMA.scala 120:63]
  wire [20:0] _T_557; // @[PositFMA.scala 121:50]
  wire [21:0] signSumSig; // @[Cat.scala 29:58]
  wire [20:0] _T_558; // @[PositFMA.scala 125:33]
  wire [20:0] _T_559; // @[PositFMA.scala 125:68]
  wire [20:0] sumXor; // @[PositFMA.scala 125:51]
  wire [15:0] _T_560; // @[LZD.scala 43:32]
  wire [7:0] _T_561; // @[LZD.scala 43:32]
  wire [3:0] _T_562; // @[LZD.scala 43:32]
  wire [1:0] _T_563; // @[LZD.scala 43:32]
  wire  _T_564; // @[LZD.scala 39:14]
  wire  _T_565; // @[LZD.scala 39:21]
  wire  _T_566; // @[LZD.scala 39:30]
  wire  _T_567; // @[LZD.scala 39:27]
  wire  _T_568; // @[LZD.scala 39:25]
  wire [1:0] _T_569; // @[Cat.scala 29:58]
  wire [1:0] _T_570; // @[LZD.scala 44:32]
  wire  _T_571; // @[LZD.scala 39:14]
  wire  _T_572; // @[LZD.scala 39:21]
  wire  _T_573; // @[LZD.scala 39:30]
  wire  _T_574; // @[LZD.scala 39:27]
  wire  _T_575; // @[LZD.scala 39:25]
  wire [1:0] _T_576; // @[Cat.scala 29:58]
  wire  _T_577; // @[Shift.scala 12:21]
  wire  _T_578; // @[Shift.scala 12:21]
  wire  _T_579; // @[LZD.scala 49:16]
  wire  _T_580; // @[LZD.scala 49:27]
  wire  _T_581; // @[LZD.scala 49:25]
  wire  _T_582; // @[LZD.scala 49:47]
  wire  _T_583; // @[LZD.scala 49:59]
  wire  _T_584; // @[LZD.scala 49:35]
  wire [2:0] _T_586; // @[Cat.scala 29:58]
  wire [3:0] _T_587; // @[LZD.scala 44:32]
  wire [1:0] _T_588; // @[LZD.scala 43:32]
  wire  _T_589; // @[LZD.scala 39:14]
  wire  _T_590; // @[LZD.scala 39:21]
  wire  _T_591; // @[LZD.scala 39:30]
  wire  _T_592; // @[LZD.scala 39:27]
  wire  _T_593; // @[LZD.scala 39:25]
  wire [1:0] _T_594; // @[Cat.scala 29:58]
  wire [1:0] _T_595; // @[LZD.scala 44:32]
  wire  _T_596; // @[LZD.scala 39:14]
  wire  _T_597; // @[LZD.scala 39:21]
  wire  _T_598; // @[LZD.scala 39:30]
  wire  _T_599; // @[LZD.scala 39:27]
  wire  _T_600; // @[LZD.scala 39:25]
  wire [1:0] _T_601; // @[Cat.scala 29:58]
  wire  _T_602; // @[Shift.scala 12:21]
  wire  _T_603; // @[Shift.scala 12:21]
  wire  _T_604; // @[LZD.scala 49:16]
  wire  _T_605; // @[LZD.scala 49:27]
  wire  _T_606; // @[LZD.scala 49:25]
  wire  _T_607; // @[LZD.scala 49:47]
  wire  _T_608; // @[LZD.scala 49:59]
  wire  _T_609; // @[LZD.scala 49:35]
  wire [2:0] _T_611; // @[Cat.scala 29:58]
  wire  _T_612; // @[Shift.scala 12:21]
  wire  _T_613; // @[Shift.scala 12:21]
  wire  _T_614; // @[LZD.scala 49:16]
  wire  _T_615; // @[LZD.scala 49:27]
  wire  _T_616; // @[LZD.scala 49:25]
  wire [1:0] _T_617; // @[LZD.scala 49:47]
  wire [1:0] _T_618; // @[LZD.scala 49:59]
  wire [1:0] _T_619; // @[LZD.scala 49:35]
  wire [3:0] _T_621; // @[Cat.scala 29:58]
  wire [7:0] _T_622; // @[LZD.scala 44:32]
  wire [3:0] _T_623; // @[LZD.scala 43:32]
  wire [1:0] _T_624; // @[LZD.scala 43:32]
  wire  _T_625; // @[LZD.scala 39:14]
  wire  _T_626; // @[LZD.scala 39:21]
  wire  _T_627; // @[LZD.scala 39:30]
  wire  _T_628; // @[LZD.scala 39:27]
  wire  _T_629; // @[LZD.scala 39:25]
  wire [1:0] _T_630; // @[Cat.scala 29:58]
  wire [1:0] _T_631; // @[LZD.scala 44:32]
  wire  _T_632; // @[LZD.scala 39:14]
  wire  _T_633; // @[LZD.scala 39:21]
  wire  _T_634; // @[LZD.scala 39:30]
  wire  _T_635; // @[LZD.scala 39:27]
  wire  _T_636; // @[LZD.scala 39:25]
  wire [1:0] _T_637; // @[Cat.scala 29:58]
  wire  _T_638; // @[Shift.scala 12:21]
  wire  _T_639; // @[Shift.scala 12:21]
  wire  _T_640; // @[LZD.scala 49:16]
  wire  _T_641; // @[LZD.scala 49:27]
  wire  _T_642; // @[LZD.scala 49:25]
  wire  _T_643; // @[LZD.scala 49:47]
  wire  _T_644; // @[LZD.scala 49:59]
  wire  _T_645; // @[LZD.scala 49:35]
  wire [2:0] _T_647; // @[Cat.scala 29:58]
  wire [3:0] _T_648; // @[LZD.scala 44:32]
  wire [1:0] _T_649; // @[LZD.scala 43:32]
  wire  _T_650; // @[LZD.scala 39:14]
  wire  _T_651; // @[LZD.scala 39:21]
  wire  _T_652; // @[LZD.scala 39:30]
  wire  _T_653; // @[LZD.scala 39:27]
  wire  _T_654; // @[LZD.scala 39:25]
  wire [1:0] _T_655; // @[Cat.scala 29:58]
  wire [1:0] _T_656; // @[LZD.scala 44:32]
  wire  _T_657; // @[LZD.scala 39:14]
  wire  _T_658; // @[LZD.scala 39:21]
  wire  _T_659; // @[LZD.scala 39:30]
  wire  _T_660; // @[LZD.scala 39:27]
  wire  _T_661; // @[LZD.scala 39:25]
  wire [1:0] _T_662; // @[Cat.scala 29:58]
  wire  _T_663; // @[Shift.scala 12:21]
  wire  _T_664; // @[Shift.scala 12:21]
  wire  _T_665; // @[LZD.scala 49:16]
  wire  _T_666; // @[LZD.scala 49:27]
  wire  _T_667; // @[LZD.scala 49:25]
  wire  _T_668; // @[LZD.scala 49:47]
  wire  _T_669; // @[LZD.scala 49:59]
  wire  _T_670; // @[LZD.scala 49:35]
  wire [2:0] _T_672; // @[Cat.scala 29:58]
  wire  _T_673; // @[Shift.scala 12:21]
  wire  _T_674; // @[Shift.scala 12:21]
  wire  _T_675; // @[LZD.scala 49:16]
  wire  _T_676; // @[LZD.scala 49:27]
  wire  _T_677; // @[LZD.scala 49:25]
  wire [1:0] _T_678; // @[LZD.scala 49:47]
  wire [1:0] _T_679; // @[LZD.scala 49:59]
  wire [1:0] _T_680; // @[LZD.scala 49:35]
  wire [3:0] _T_682; // @[Cat.scala 29:58]
  wire  _T_683; // @[Shift.scala 12:21]
  wire  _T_684; // @[Shift.scala 12:21]
  wire  _T_685; // @[LZD.scala 49:16]
  wire  _T_686; // @[LZD.scala 49:27]
  wire  _T_687; // @[LZD.scala 49:25]
  wire [2:0] _T_688; // @[LZD.scala 49:47]
  wire [2:0] _T_689; // @[LZD.scala 49:59]
  wire [2:0] _T_690; // @[LZD.scala 49:35]
  wire [4:0] _T_692; // @[Cat.scala 29:58]
  wire [4:0] _T_693; // @[LZD.scala 44:32]
  wire [3:0] _T_694; // @[LZD.scala 43:32]
  wire [1:0] _T_695; // @[LZD.scala 43:32]
  wire  _T_696; // @[LZD.scala 39:14]
  wire  _T_697; // @[LZD.scala 39:21]
  wire  _T_698; // @[LZD.scala 39:30]
  wire  _T_699; // @[LZD.scala 39:27]
  wire  _T_700; // @[LZD.scala 39:25]
  wire [1:0] _T_701; // @[Cat.scala 29:58]
  wire [1:0] _T_702; // @[LZD.scala 44:32]
  wire  _T_703; // @[LZD.scala 39:14]
  wire  _T_704; // @[LZD.scala 39:21]
  wire  _T_705; // @[LZD.scala 39:30]
  wire  _T_706; // @[LZD.scala 39:27]
  wire  _T_707; // @[LZD.scala 39:25]
  wire [1:0] _T_708; // @[Cat.scala 29:58]
  wire  _T_709; // @[Shift.scala 12:21]
  wire  _T_710; // @[Shift.scala 12:21]
  wire  _T_711; // @[LZD.scala 49:16]
  wire  _T_712; // @[LZD.scala 49:27]
  wire  _T_713; // @[LZD.scala 49:25]
  wire  _T_714; // @[LZD.scala 49:47]
  wire  _T_715; // @[LZD.scala 49:59]
  wire  _T_716; // @[LZD.scala 49:35]
  wire [2:0] _T_718; // @[Cat.scala 29:58]
  wire  _T_719; // @[LZD.scala 44:32]
  wire  _T_721; // @[Shift.scala 12:21]
  wire [1:0] _T_723; // @[Cat.scala 29:58]
  wire [1:0] _T_724; // @[LZD.scala 55:32]
  wire [1:0] _T_725; // @[LZD.scala 55:20]
  wire  _T_727; // @[Shift.scala 12:21]
  wire [3:0] _T_729; // @[Cat.scala 29:58]
  wire [3:0] _T_730; // @[LZD.scala 55:32]
  wire [3:0] _T_731; // @[LZD.scala 55:20]
  wire [4:0] sumLZD; // @[Cat.scala 29:58]
  wire [4:0] shiftValue; // @[PositFMA.scala 127:24]
  wire [19:0] _T_732; // @[PositFMA.scala 128:38]
  wire  _T_733; // @[Shift.scala 16:24]
  wire  _T_735; // @[Shift.scala 12:21]
  wire [3:0] _T_736; // @[Shift.scala 64:52]
  wire [19:0] _T_738; // @[Cat.scala 29:58]
  wire [19:0] _T_739; // @[Shift.scala 64:27]
  wire [3:0] _T_740; // @[Shift.scala 66:70]
  wire  _T_741; // @[Shift.scala 12:21]
  wire [11:0] _T_742; // @[Shift.scala 64:52]
  wire [19:0] _T_744; // @[Cat.scala 29:58]
  wire [19:0] _T_745; // @[Shift.scala 64:27]
  wire [2:0] _T_746; // @[Shift.scala 66:70]
  wire  _T_747; // @[Shift.scala 12:21]
  wire [15:0] _T_748; // @[Shift.scala 64:52]
  wire [19:0] _T_750; // @[Cat.scala 29:58]
  wire [19:0] _T_751; // @[Shift.scala 64:27]
  wire [1:0] _T_752; // @[Shift.scala 66:70]
  wire  _T_753; // @[Shift.scala 12:21]
  wire [17:0] _T_754; // @[Shift.scala 64:52]
  wire [19:0] _T_756; // @[Cat.scala 29:58]
  wire [19:0] _T_757; // @[Shift.scala 64:27]
  wire  _T_758; // @[Shift.scala 66:70]
  wire [18:0] _T_760; // @[Shift.scala 64:52]
  wire [19:0] _T_761; // @[Cat.scala 29:58]
  wire [19:0] _T_762; // @[Shift.scala 64:27]
  wire [19:0] normalFracTmp; // @[Shift.scala 16:10]
  wire [6:0] _T_764; // @[PositFMA.scala 131:36]
  wire [6:0] _T_765; // @[PositFMA.scala 131:36]
  wire [5:0] _T_766; // @[Cat.scala 29:58]
  wire [5:0] _T_767; // @[PositFMA.scala 131:61]
  wire [6:0] _GEN_19; // @[PositFMA.scala 131:42]
  wire [6:0] _T_769; // @[PositFMA.scala 131:42]
  wire [6:0] sumScale; // @[PositFMA.scala 131:42]
  wire [8:0] sumFrac; // @[PositFMA.scala 132:41]
  wire [10:0] grsTmp; // @[PositFMA.scala 135:41]
  wire [1:0] _T_770; // @[PositFMA.scala 138:40]
  wire [8:0] _T_771; // @[PositFMA.scala 138:56]
  wire  _T_772; // @[PositFMA.scala 138:60]
  wire  underflow; // @[PositFMA.scala 145:32]
  wire  overflow; // @[PositFMA.scala 146:32]
  wire  _T_773; // @[PositFMA.scala 155:32]
  wire  decF_isZero; // @[PositFMA.scala 155:20]
  wire [6:0] _T_775; // @[Mux.scala 87:16]
  wire [6:0] _T_776; // @[Mux.scala 87:16]
  wire [5:0] _GEN_20; // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  wire [5:0] decF_scale; // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  wire  _T_777; // @[convert.scala 46:61]
  wire  _T_778; // @[convert.scala 46:52]
  wire  _T_780; // @[convert.scala 46:42]
  wire [4:0] _T_781; // @[convert.scala 48:34]
  wire  _T_782; // @[convert.scala 49:36]
  wire [4:0] _T_784; // @[convert.scala 50:36]
  wire [4:0] _T_785; // @[convert.scala 50:36]
  wire [4:0] _T_786; // @[convert.scala 50:28]
  wire  _T_787; // @[convert.scala 51:31]
  wire  _T_788; // @[convert.scala 52:43]
  wire [14:0] _T_792; // @[Cat.scala 29:58]
  wire [4:0] _T_793; // @[Shift.scala 39:17]
  wire  _T_794; // @[Shift.scala 39:24]
  wire [3:0] _T_795; // @[Shift.scala 40:44]
  wire [6:0] _T_796; // @[Shift.scala 90:30]
  wire [7:0] _T_797; // @[Shift.scala 90:48]
  wire  _T_798; // @[Shift.scala 90:57]
  wire [6:0] _GEN_21; // @[Shift.scala 90:39]
  wire [6:0] _T_799; // @[Shift.scala 90:39]
  wire  _T_800; // @[Shift.scala 12:21]
  wire  _T_801; // @[Shift.scala 12:21]
  wire [7:0] _T_803; // @[Bitwise.scala 71:12]
  wire [14:0] _T_804; // @[Cat.scala 29:58]
  wire [14:0] _T_805; // @[Shift.scala 91:22]
  wire [2:0] _T_806; // @[Shift.scala 92:77]
  wire [10:0] _T_807; // @[Shift.scala 90:30]
  wire [3:0] _T_808; // @[Shift.scala 90:48]
  wire  _T_809; // @[Shift.scala 90:57]
  wire [10:0] _GEN_22; // @[Shift.scala 90:39]
  wire [10:0] _T_810; // @[Shift.scala 90:39]
  wire  _T_811; // @[Shift.scala 12:21]
  wire  _T_812; // @[Shift.scala 12:21]
  wire [3:0] _T_814; // @[Bitwise.scala 71:12]
  wire [14:0] _T_815; // @[Cat.scala 29:58]
  wire [14:0] _T_816; // @[Shift.scala 91:22]
  wire [1:0] _T_817; // @[Shift.scala 92:77]
  wire [12:0] _T_818; // @[Shift.scala 90:30]
  wire [1:0] _T_819; // @[Shift.scala 90:48]
  wire  _T_820; // @[Shift.scala 90:57]
  wire [12:0] _GEN_23; // @[Shift.scala 90:39]
  wire [12:0] _T_821; // @[Shift.scala 90:39]
  wire  _T_822; // @[Shift.scala 12:21]
  wire  _T_823; // @[Shift.scala 12:21]
  wire [1:0] _T_825; // @[Bitwise.scala 71:12]
  wire [14:0] _T_826; // @[Cat.scala 29:58]
  wire [14:0] _T_827; // @[Shift.scala 91:22]
  wire  _T_828; // @[Shift.scala 92:77]
  wire [13:0] _T_829; // @[Shift.scala 90:30]
  wire  _T_830; // @[Shift.scala 90:48]
  wire [13:0] _GEN_24; // @[Shift.scala 90:39]
  wire [13:0] _T_832; // @[Shift.scala 90:39]
  wire  _T_834; // @[Shift.scala 12:21]
  wire [14:0] _T_835; // @[Cat.scala 29:58]
  wire [14:0] _T_836; // @[Shift.scala 91:22]
  wire [14:0] _T_839; // @[Bitwise.scala 71:12]
  wire [14:0] _T_840; // @[Shift.scala 39:10]
  wire  _T_841; // @[convert.scala 55:31]
  wire  _T_842; // @[convert.scala 56:31]
  wire  _T_843; // @[convert.scala 57:31]
  wire  _T_844; // @[convert.scala 58:31]
  wire [11:0] _T_845; // @[convert.scala 59:69]
  wire  _T_846; // @[convert.scala 59:81]
  wire  _T_847; // @[convert.scala 59:50]
  wire  _T_849; // @[convert.scala 60:81]
  wire  _T_850; // @[convert.scala 61:44]
  wire  _T_851; // @[convert.scala 61:52]
  wire  _T_852; // @[convert.scala 61:36]
  wire  _T_853; // @[convert.scala 62:63]
  wire  _T_854; // @[convert.scala 62:103]
  wire  _T_855; // @[convert.scala 62:60]
  wire [11:0] _GEN_25; // @[convert.scala 63:56]
  wire [11:0] _T_858; // @[convert.scala 63:56]
  wire [12:0] _T_859; // @[Cat.scala 29:58]
  reg  _T_863; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [12:0] _T_867; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  assign _T = io_fmaOp[1]; // @[PositFMA.scala 47:36]
  assign _T_2 = _T ? 13'h1fff : 13'h0; // @[Bitwise.scala 71:12]
  assign _T_3 = _T_2 ^ io_A; // @[PositFMA.scala 47:41]
  assign _GEN_10 = {{12'd0}, _T}; // @[PositFMA.scala 47:49]
  assign realA = _T_3 + _GEN_10; // @[PositFMA.scala 47:49]
  assign _T_6 = io_fmaOp[0]; // @[PositFMA.scala 48:36]
  assign _T_8 = _T_6 ? 13'h1fff : 13'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = _T_8 ^ io_C; // @[PositFMA.scala 48:41]
  assign _GEN_11 = {{12'd0}, _T_6}; // @[PositFMA.scala 48:49]
  assign realC = _T_9 + _GEN_11; // @[PositFMA.scala 48:49]
  assign _T_13 = realA[12]; // @[convert.scala 18:24]
  assign _T_14 = realA[11]; // @[convert.scala 18:40]
  assign _T_15 = _T_13 ^ _T_14; // @[convert.scala 18:36]
  assign _T_16 = realA[11:1]; // @[convert.scala 19:24]
  assign _T_17 = realA[10:0]; // @[convert.scala 19:43]
  assign _T_18 = _T_16 ^ _T_17; // @[convert.scala 19:39]
  assign _T_19 = _T_18[10:3]; // @[LZD.scala 43:32]
  assign _T_20 = _T_19[7:4]; // @[LZD.scala 43:32]
  assign _T_21 = _T_20[3:2]; // @[LZD.scala 43:32]
  assign _T_22 = _T_21 != 2'h0; // @[LZD.scala 39:14]
  assign _T_23 = _T_21[1]; // @[LZD.scala 39:21]
  assign _T_24 = _T_21[0]; // @[LZD.scala 39:30]
  assign _T_25 = ~ _T_24; // @[LZD.scala 39:27]
  assign _T_26 = _T_23 | _T_25; // @[LZD.scala 39:25]
  assign _T_27 = {_T_22,_T_26}; // @[Cat.scala 29:58]
  assign _T_28 = _T_20[1:0]; // @[LZD.scala 44:32]
  assign _T_29 = _T_28 != 2'h0; // @[LZD.scala 39:14]
  assign _T_30 = _T_28[1]; // @[LZD.scala 39:21]
  assign _T_31 = _T_28[0]; // @[LZD.scala 39:30]
  assign _T_32 = ~ _T_31; // @[LZD.scala 39:27]
  assign _T_33 = _T_30 | _T_32; // @[LZD.scala 39:25]
  assign _T_34 = {_T_29,_T_33}; // @[Cat.scala 29:58]
  assign _T_35 = _T_27[1]; // @[Shift.scala 12:21]
  assign _T_36 = _T_34[1]; // @[Shift.scala 12:21]
  assign _T_37 = _T_35 | _T_36; // @[LZD.scala 49:16]
  assign _T_38 = ~ _T_36; // @[LZD.scala 49:27]
  assign _T_39 = _T_35 | _T_38; // @[LZD.scala 49:25]
  assign _T_40 = _T_27[0:0]; // @[LZD.scala 49:47]
  assign _T_41 = _T_34[0:0]; // @[LZD.scala 49:59]
  assign _T_42 = _T_35 ? _T_40 : _T_41; // @[LZD.scala 49:35]
  assign _T_44 = {_T_37,_T_39,_T_42}; // @[Cat.scala 29:58]
  assign _T_45 = _T_19[3:0]; // @[LZD.scala 44:32]
  assign _T_46 = _T_45[3:2]; // @[LZD.scala 43:32]
  assign _T_47 = _T_46 != 2'h0; // @[LZD.scala 39:14]
  assign _T_48 = _T_46[1]; // @[LZD.scala 39:21]
  assign _T_49 = _T_46[0]; // @[LZD.scala 39:30]
  assign _T_50 = ~ _T_49; // @[LZD.scala 39:27]
  assign _T_51 = _T_48 | _T_50; // @[LZD.scala 39:25]
  assign _T_52 = {_T_47,_T_51}; // @[Cat.scala 29:58]
  assign _T_53 = _T_45[1:0]; // @[LZD.scala 44:32]
  assign _T_54 = _T_53 != 2'h0; // @[LZD.scala 39:14]
  assign _T_55 = _T_53[1]; // @[LZD.scala 39:21]
  assign _T_56 = _T_53[0]; // @[LZD.scala 39:30]
  assign _T_57 = ~ _T_56; // @[LZD.scala 39:27]
  assign _T_58 = _T_55 | _T_57; // @[LZD.scala 39:25]
  assign _T_59 = {_T_54,_T_58}; // @[Cat.scala 29:58]
  assign _T_60 = _T_52[1]; // @[Shift.scala 12:21]
  assign _T_61 = _T_59[1]; // @[Shift.scala 12:21]
  assign _T_62 = _T_60 | _T_61; // @[LZD.scala 49:16]
  assign _T_63 = ~ _T_61; // @[LZD.scala 49:27]
  assign _T_64 = _T_60 | _T_63; // @[LZD.scala 49:25]
  assign _T_65 = _T_52[0:0]; // @[LZD.scala 49:47]
  assign _T_66 = _T_59[0:0]; // @[LZD.scala 49:59]
  assign _T_67 = _T_60 ? _T_65 : _T_66; // @[LZD.scala 49:35]
  assign _T_69 = {_T_62,_T_64,_T_67}; // @[Cat.scala 29:58]
  assign _T_70 = _T_44[2]; // @[Shift.scala 12:21]
  assign _T_71 = _T_69[2]; // @[Shift.scala 12:21]
  assign _T_72 = _T_70 | _T_71; // @[LZD.scala 49:16]
  assign _T_73 = ~ _T_71; // @[LZD.scala 49:27]
  assign _T_74 = _T_70 | _T_73; // @[LZD.scala 49:25]
  assign _T_75 = _T_44[1:0]; // @[LZD.scala 49:47]
  assign _T_76 = _T_69[1:0]; // @[LZD.scala 49:59]
  assign _T_77 = _T_70 ? _T_75 : _T_76; // @[LZD.scala 49:35]
  assign _T_79 = {_T_72,_T_74,_T_77}; // @[Cat.scala 29:58]
  assign _T_80 = _T_18[2:0]; // @[LZD.scala 44:32]
  assign _T_81 = _T_80[2:1]; // @[LZD.scala 43:32]
  assign _T_82 = _T_81 != 2'h0; // @[LZD.scala 39:14]
  assign _T_83 = _T_81[1]; // @[LZD.scala 39:21]
  assign _T_84 = _T_81[0]; // @[LZD.scala 39:30]
  assign _T_85 = ~ _T_84; // @[LZD.scala 39:27]
  assign _T_86 = _T_83 | _T_85; // @[LZD.scala 39:25]
  assign _T_87 = {_T_82,_T_86}; // @[Cat.scala 29:58]
  assign _T_88 = _T_80[0:0]; // @[LZD.scala 44:32]
  assign _T_90 = _T_87[1]; // @[Shift.scala 12:21]
  assign _T_92 = _T_87[0:0]; // @[LZD.scala 55:32]
  assign _T_93 = _T_90 ? _T_92 : _T_88; // @[LZD.scala 55:20]
  assign _T_95 = _T_79[3]; // @[Shift.scala 12:21]
  assign _T_97 = {1'h1,_T_90,_T_93}; // @[Cat.scala 29:58]
  assign _T_98 = _T_79[2:0]; // @[LZD.scala 55:32]
  assign _T_99 = _T_95 ? _T_98 : _T_97; // @[LZD.scala 55:20]
  assign _T_100 = {_T_95,_T_99}; // @[Cat.scala 29:58]
  assign _T_101 = ~ _T_100; // @[convert.scala 21:22]
  assign _T_102 = realA[9:0]; // @[convert.scala 22:36]
  assign _T_103 = _T_101 < 4'ha; // @[Shift.scala 16:24]
  assign _T_105 = _T_101[3]; // @[Shift.scala 12:21]
  assign _T_106 = _T_102[1:0]; // @[Shift.scala 64:52]
  assign _T_108 = {_T_106,8'h0}; // @[Cat.scala 29:58]
  assign _T_109 = _T_105 ? _T_108 : _T_102; // @[Shift.scala 64:27]
  assign _T_110 = _T_101[2:0]; // @[Shift.scala 66:70]
  assign _T_111 = _T_110[2]; // @[Shift.scala 12:21]
  assign _T_112 = _T_109[5:0]; // @[Shift.scala 64:52]
  assign _T_114 = {_T_112,4'h0}; // @[Cat.scala 29:58]
  assign _T_115 = _T_111 ? _T_114 : _T_109; // @[Shift.scala 64:27]
  assign _T_116 = _T_110[1:0]; // @[Shift.scala 66:70]
  assign _T_117 = _T_116[1]; // @[Shift.scala 12:21]
  assign _T_118 = _T_115[7:0]; // @[Shift.scala 64:52]
  assign _T_120 = {_T_118,2'h0}; // @[Cat.scala 29:58]
  assign _T_121 = _T_117 ? _T_120 : _T_115; // @[Shift.scala 64:27]
  assign _T_122 = _T_116[0:0]; // @[Shift.scala 66:70]
  assign _T_124 = _T_121[8:0]; // @[Shift.scala 64:52]
  assign _T_125 = {_T_124,1'h0}; // @[Cat.scala 29:58]
  assign _T_126 = _T_122 ? _T_125 : _T_121; // @[Shift.scala 64:27]
  assign _T_127 = _T_103 ? _T_126 : 10'h0; // @[Shift.scala 16:10]
  assign _T_128 = _T_127[9:9]; // @[convert.scala 23:34]
  assign decA_fraction = _T_127[8:0]; // @[convert.scala 24:34]
  assign _T_130 = _T_15 == 1'h0; // @[convert.scala 25:26]
  assign _T_132 = _T_15 ? _T_101 : _T_100; // @[convert.scala 25:42]
  assign _T_135 = ~ _T_128; // @[convert.scala 26:67]
  assign _T_136 = _T_13 ? _T_135 : _T_128; // @[convert.scala 26:51]
  assign _T_137 = {_T_130,_T_132,_T_136}; // @[Cat.scala 29:58]
  assign _T_139 = realA[11:0]; // @[convert.scala 29:56]
  assign _T_140 = _T_139 != 12'h0; // @[convert.scala 29:60]
  assign _T_141 = ~ _T_140; // @[convert.scala 29:41]
  assign decA_isNaR = _T_13 & _T_141; // @[convert.scala 29:39]
  assign _T_144 = _T_13 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_144 & _T_141; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_137); // @[convert.scala 32:24]
  assign _T_153 = io_B[12]; // @[convert.scala 18:24]
  assign _T_154 = io_B[11]; // @[convert.scala 18:40]
  assign _T_155 = _T_153 ^ _T_154; // @[convert.scala 18:36]
  assign _T_156 = io_B[11:1]; // @[convert.scala 19:24]
  assign _T_157 = io_B[10:0]; // @[convert.scala 19:43]
  assign _T_158 = _T_156 ^ _T_157; // @[convert.scala 19:39]
  assign _T_159 = _T_158[10:3]; // @[LZD.scala 43:32]
  assign _T_160 = _T_159[7:4]; // @[LZD.scala 43:32]
  assign _T_161 = _T_160[3:2]; // @[LZD.scala 43:32]
  assign _T_162 = _T_161 != 2'h0; // @[LZD.scala 39:14]
  assign _T_163 = _T_161[1]; // @[LZD.scala 39:21]
  assign _T_164 = _T_161[0]; // @[LZD.scala 39:30]
  assign _T_165 = ~ _T_164; // @[LZD.scala 39:27]
  assign _T_166 = _T_163 | _T_165; // @[LZD.scala 39:25]
  assign _T_167 = {_T_162,_T_166}; // @[Cat.scala 29:58]
  assign _T_168 = _T_160[1:0]; // @[LZD.scala 44:32]
  assign _T_169 = _T_168 != 2'h0; // @[LZD.scala 39:14]
  assign _T_170 = _T_168[1]; // @[LZD.scala 39:21]
  assign _T_171 = _T_168[0]; // @[LZD.scala 39:30]
  assign _T_172 = ~ _T_171; // @[LZD.scala 39:27]
  assign _T_173 = _T_170 | _T_172; // @[LZD.scala 39:25]
  assign _T_174 = {_T_169,_T_173}; // @[Cat.scala 29:58]
  assign _T_175 = _T_167[1]; // @[Shift.scala 12:21]
  assign _T_176 = _T_174[1]; // @[Shift.scala 12:21]
  assign _T_177 = _T_175 | _T_176; // @[LZD.scala 49:16]
  assign _T_178 = ~ _T_176; // @[LZD.scala 49:27]
  assign _T_179 = _T_175 | _T_178; // @[LZD.scala 49:25]
  assign _T_180 = _T_167[0:0]; // @[LZD.scala 49:47]
  assign _T_181 = _T_174[0:0]; // @[LZD.scala 49:59]
  assign _T_182 = _T_175 ? _T_180 : _T_181; // @[LZD.scala 49:35]
  assign _T_184 = {_T_177,_T_179,_T_182}; // @[Cat.scala 29:58]
  assign _T_185 = _T_159[3:0]; // @[LZD.scala 44:32]
  assign _T_186 = _T_185[3:2]; // @[LZD.scala 43:32]
  assign _T_187 = _T_186 != 2'h0; // @[LZD.scala 39:14]
  assign _T_188 = _T_186[1]; // @[LZD.scala 39:21]
  assign _T_189 = _T_186[0]; // @[LZD.scala 39:30]
  assign _T_190 = ~ _T_189; // @[LZD.scala 39:27]
  assign _T_191 = _T_188 | _T_190; // @[LZD.scala 39:25]
  assign _T_192 = {_T_187,_T_191}; // @[Cat.scala 29:58]
  assign _T_193 = _T_185[1:0]; // @[LZD.scala 44:32]
  assign _T_194 = _T_193 != 2'h0; // @[LZD.scala 39:14]
  assign _T_195 = _T_193[1]; // @[LZD.scala 39:21]
  assign _T_196 = _T_193[0]; // @[LZD.scala 39:30]
  assign _T_197 = ~ _T_196; // @[LZD.scala 39:27]
  assign _T_198 = _T_195 | _T_197; // @[LZD.scala 39:25]
  assign _T_199 = {_T_194,_T_198}; // @[Cat.scala 29:58]
  assign _T_200 = _T_192[1]; // @[Shift.scala 12:21]
  assign _T_201 = _T_199[1]; // @[Shift.scala 12:21]
  assign _T_202 = _T_200 | _T_201; // @[LZD.scala 49:16]
  assign _T_203 = ~ _T_201; // @[LZD.scala 49:27]
  assign _T_204 = _T_200 | _T_203; // @[LZD.scala 49:25]
  assign _T_205 = _T_192[0:0]; // @[LZD.scala 49:47]
  assign _T_206 = _T_199[0:0]; // @[LZD.scala 49:59]
  assign _T_207 = _T_200 ? _T_205 : _T_206; // @[LZD.scala 49:35]
  assign _T_209 = {_T_202,_T_204,_T_207}; // @[Cat.scala 29:58]
  assign _T_210 = _T_184[2]; // @[Shift.scala 12:21]
  assign _T_211 = _T_209[2]; // @[Shift.scala 12:21]
  assign _T_212 = _T_210 | _T_211; // @[LZD.scala 49:16]
  assign _T_213 = ~ _T_211; // @[LZD.scala 49:27]
  assign _T_214 = _T_210 | _T_213; // @[LZD.scala 49:25]
  assign _T_215 = _T_184[1:0]; // @[LZD.scala 49:47]
  assign _T_216 = _T_209[1:0]; // @[LZD.scala 49:59]
  assign _T_217 = _T_210 ? _T_215 : _T_216; // @[LZD.scala 49:35]
  assign _T_219 = {_T_212,_T_214,_T_217}; // @[Cat.scala 29:58]
  assign _T_220 = _T_158[2:0]; // @[LZD.scala 44:32]
  assign _T_221 = _T_220[2:1]; // @[LZD.scala 43:32]
  assign _T_222 = _T_221 != 2'h0; // @[LZD.scala 39:14]
  assign _T_223 = _T_221[1]; // @[LZD.scala 39:21]
  assign _T_224 = _T_221[0]; // @[LZD.scala 39:30]
  assign _T_225 = ~ _T_224; // @[LZD.scala 39:27]
  assign _T_226 = _T_223 | _T_225; // @[LZD.scala 39:25]
  assign _T_227 = {_T_222,_T_226}; // @[Cat.scala 29:58]
  assign _T_228 = _T_220[0:0]; // @[LZD.scala 44:32]
  assign _T_230 = _T_227[1]; // @[Shift.scala 12:21]
  assign _T_232 = _T_227[0:0]; // @[LZD.scala 55:32]
  assign _T_233 = _T_230 ? _T_232 : _T_228; // @[LZD.scala 55:20]
  assign _T_235 = _T_219[3]; // @[Shift.scala 12:21]
  assign _T_237 = {1'h1,_T_230,_T_233}; // @[Cat.scala 29:58]
  assign _T_238 = _T_219[2:0]; // @[LZD.scala 55:32]
  assign _T_239 = _T_235 ? _T_238 : _T_237; // @[LZD.scala 55:20]
  assign _T_240 = {_T_235,_T_239}; // @[Cat.scala 29:58]
  assign _T_241 = ~ _T_240; // @[convert.scala 21:22]
  assign _T_242 = io_B[9:0]; // @[convert.scala 22:36]
  assign _T_243 = _T_241 < 4'ha; // @[Shift.scala 16:24]
  assign _T_245 = _T_241[3]; // @[Shift.scala 12:21]
  assign _T_246 = _T_242[1:0]; // @[Shift.scala 64:52]
  assign _T_248 = {_T_246,8'h0}; // @[Cat.scala 29:58]
  assign _T_249 = _T_245 ? _T_248 : _T_242; // @[Shift.scala 64:27]
  assign _T_250 = _T_241[2:0]; // @[Shift.scala 66:70]
  assign _T_251 = _T_250[2]; // @[Shift.scala 12:21]
  assign _T_252 = _T_249[5:0]; // @[Shift.scala 64:52]
  assign _T_254 = {_T_252,4'h0}; // @[Cat.scala 29:58]
  assign _T_255 = _T_251 ? _T_254 : _T_249; // @[Shift.scala 64:27]
  assign _T_256 = _T_250[1:0]; // @[Shift.scala 66:70]
  assign _T_257 = _T_256[1]; // @[Shift.scala 12:21]
  assign _T_258 = _T_255[7:0]; // @[Shift.scala 64:52]
  assign _T_260 = {_T_258,2'h0}; // @[Cat.scala 29:58]
  assign _T_261 = _T_257 ? _T_260 : _T_255; // @[Shift.scala 64:27]
  assign _T_262 = _T_256[0:0]; // @[Shift.scala 66:70]
  assign _T_264 = _T_261[8:0]; // @[Shift.scala 64:52]
  assign _T_265 = {_T_264,1'h0}; // @[Cat.scala 29:58]
  assign _T_266 = _T_262 ? _T_265 : _T_261; // @[Shift.scala 64:27]
  assign _T_267 = _T_243 ? _T_266 : 10'h0; // @[Shift.scala 16:10]
  assign _T_268 = _T_267[9:9]; // @[convert.scala 23:34]
  assign decB_fraction = _T_267[8:0]; // @[convert.scala 24:34]
  assign _T_270 = _T_155 == 1'h0; // @[convert.scala 25:26]
  assign _T_272 = _T_155 ? _T_241 : _T_240; // @[convert.scala 25:42]
  assign _T_275 = ~ _T_268; // @[convert.scala 26:67]
  assign _T_276 = _T_153 ? _T_275 : _T_268; // @[convert.scala 26:51]
  assign _T_277 = {_T_270,_T_272,_T_276}; // @[Cat.scala 29:58]
  assign _T_279 = io_B[11:0]; // @[convert.scala 29:56]
  assign _T_280 = _T_279 != 12'h0; // @[convert.scala 29:60]
  assign _T_281 = ~ _T_280; // @[convert.scala 29:41]
  assign decB_isNaR = _T_153 & _T_281; // @[convert.scala 29:39]
  assign _T_284 = _T_153 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_284 & _T_281; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_277); // @[convert.scala 32:24]
  assign _T_293 = realC[12]; // @[convert.scala 18:24]
  assign _T_294 = realC[11]; // @[convert.scala 18:40]
  assign _T_295 = _T_293 ^ _T_294; // @[convert.scala 18:36]
  assign _T_296 = realC[11:1]; // @[convert.scala 19:24]
  assign _T_297 = realC[10:0]; // @[convert.scala 19:43]
  assign _T_298 = _T_296 ^ _T_297; // @[convert.scala 19:39]
  assign _T_299 = _T_298[10:3]; // @[LZD.scala 43:32]
  assign _T_300 = _T_299[7:4]; // @[LZD.scala 43:32]
  assign _T_301 = _T_300[3:2]; // @[LZD.scala 43:32]
  assign _T_302 = _T_301 != 2'h0; // @[LZD.scala 39:14]
  assign _T_303 = _T_301[1]; // @[LZD.scala 39:21]
  assign _T_304 = _T_301[0]; // @[LZD.scala 39:30]
  assign _T_305 = ~ _T_304; // @[LZD.scala 39:27]
  assign _T_306 = _T_303 | _T_305; // @[LZD.scala 39:25]
  assign _T_307 = {_T_302,_T_306}; // @[Cat.scala 29:58]
  assign _T_308 = _T_300[1:0]; // @[LZD.scala 44:32]
  assign _T_309 = _T_308 != 2'h0; // @[LZD.scala 39:14]
  assign _T_310 = _T_308[1]; // @[LZD.scala 39:21]
  assign _T_311 = _T_308[0]; // @[LZD.scala 39:30]
  assign _T_312 = ~ _T_311; // @[LZD.scala 39:27]
  assign _T_313 = _T_310 | _T_312; // @[LZD.scala 39:25]
  assign _T_314 = {_T_309,_T_313}; // @[Cat.scala 29:58]
  assign _T_315 = _T_307[1]; // @[Shift.scala 12:21]
  assign _T_316 = _T_314[1]; // @[Shift.scala 12:21]
  assign _T_317 = _T_315 | _T_316; // @[LZD.scala 49:16]
  assign _T_318 = ~ _T_316; // @[LZD.scala 49:27]
  assign _T_319 = _T_315 | _T_318; // @[LZD.scala 49:25]
  assign _T_320 = _T_307[0:0]; // @[LZD.scala 49:47]
  assign _T_321 = _T_314[0:0]; // @[LZD.scala 49:59]
  assign _T_322 = _T_315 ? _T_320 : _T_321; // @[LZD.scala 49:35]
  assign _T_324 = {_T_317,_T_319,_T_322}; // @[Cat.scala 29:58]
  assign _T_325 = _T_299[3:0]; // @[LZD.scala 44:32]
  assign _T_326 = _T_325[3:2]; // @[LZD.scala 43:32]
  assign _T_327 = _T_326 != 2'h0; // @[LZD.scala 39:14]
  assign _T_328 = _T_326[1]; // @[LZD.scala 39:21]
  assign _T_329 = _T_326[0]; // @[LZD.scala 39:30]
  assign _T_330 = ~ _T_329; // @[LZD.scala 39:27]
  assign _T_331 = _T_328 | _T_330; // @[LZD.scala 39:25]
  assign _T_332 = {_T_327,_T_331}; // @[Cat.scala 29:58]
  assign _T_333 = _T_325[1:0]; // @[LZD.scala 44:32]
  assign _T_334 = _T_333 != 2'h0; // @[LZD.scala 39:14]
  assign _T_335 = _T_333[1]; // @[LZD.scala 39:21]
  assign _T_336 = _T_333[0]; // @[LZD.scala 39:30]
  assign _T_337 = ~ _T_336; // @[LZD.scala 39:27]
  assign _T_338 = _T_335 | _T_337; // @[LZD.scala 39:25]
  assign _T_339 = {_T_334,_T_338}; // @[Cat.scala 29:58]
  assign _T_340 = _T_332[1]; // @[Shift.scala 12:21]
  assign _T_341 = _T_339[1]; // @[Shift.scala 12:21]
  assign _T_342 = _T_340 | _T_341; // @[LZD.scala 49:16]
  assign _T_343 = ~ _T_341; // @[LZD.scala 49:27]
  assign _T_344 = _T_340 | _T_343; // @[LZD.scala 49:25]
  assign _T_345 = _T_332[0:0]; // @[LZD.scala 49:47]
  assign _T_346 = _T_339[0:0]; // @[LZD.scala 49:59]
  assign _T_347 = _T_340 ? _T_345 : _T_346; // @[LZD.scala 49:35]
  assign _T_349 = {_T_342,_T_344,_T_347}; // @[Cat.scala 29:58]
  assign _T_350 = _T_324[2]; // @[Shift.scala 12:21]
  assign _T_351 = _T_349[2]; // @[Shift.scala 12:21]
  assign _T_352 = _T_350 | _T_351; // @[LZD.scala 49:16]
  assign _T_353 = ~ _T_351; // @[LZD.scala 49:27]
  assign _T_354 = _T_350 | _T_353; // @[LZD.scala 49:25]
  assign _T_355 = _T_324[1:0]; // @[LZD.scala 49:47]
  assign _T_356 = _T_349[1:0]; // @[LZD.scala 49:59]
  assign _T_357 = _T_350 ? _T_355 : _T_356; // @[LZD.scala 49:35]
  assign _T_359 = {_T_352,_T_354,_T_357}; // @[Cat.scala 29:58]
  assign _T_360 = _T_298[2:0]; // @[LZD.scala 44:32]
  assign _T_361 = _T_360[2:1]; // @[LZD.scala 43:32]
  assign _T_362 = _T_361 != 2'h0; // @[LZD.scala 39:14]
  assign _T_363 = _T_361[1]; // @[LZD.scala 39:21]
  assign _T_364 = _T_361[0]; // @[LZD.scala 39:30]
  assign _T_365 = ~ _T_364; // @[LZD.scala 39:27]
  assign _T_366 = _T_363 | _T_365; // @[LZD.scala 39:25]
  assign _T_367 = {_T_362,_T_366}; // @[Cat.scala 29:58]
  assign _T_368 = _T_360[0:0]; // @[LZD.scala 44:32]
  assign _T_370 = _T_367[1]; // @[Shift.scala 12:21]
  assign _T_372 = _T_367[0:0]; // @[LZD.scala 55:32]
  assign _T_373 = _T_370 ? _T_372 : _T_368; // @[LZD.scala 55:20]
  assign _T_375 = _T_359[3]; // @[Shift.scala 12:21]
  assign _T_377 = {1'h1,_T_370,_T_373}; // @[Cat.scala 29:58]
  assign _T_378 = _T_359[2:0]; // @[LZD.scala 55:32]
  assign _T_379 = _T_375 ? _T_378 : _T_377; // @[LZD.scala 55:20]
  assign _T_380 = {_T_375,_T_379}; // @[Cat.scala 29:58]
  assign _T_381 = ~ _T_380; // @[convert.scala 21:22]
  assign _T_382 = realC[9:0]; // @[convert.scala 22:36]
  assign _T_383 = _T_381 < 4'ha; // @[Shift.scala 16:24]
  assign _T_385 = _T_381[3]; // @[Shift.scala 12:21]
  assign _T_386 = _T_382[1:0]; // @[Shift.scala 64:52]
  assign _T_388 = {_T_386,8'h0}; // @[Cat.scala 29:58]
  assign _T_389 = _T_385 ? _T_388 : _T_382; // @[Shift.scala 64:27]
  assign _T_390 = _T_381[2:0]; // @[Shift.scala 66:70]
  assign _T_391 = _T_390[2]; // @[Shift.scala 12:21]
  assign _T_392 = _T_389[5:0]; // @[Shift.scala 64:52]
  assign _T_394 = {_T_392,4'h0}; // @[Cat.scala 29:58]
  assign _T_395 = _T_391 ? _T_394 : _T_389; // @[Shift.scala 64:27]
  assign _T_396 = _T_390[1:0]; // @[Shift.scala 66:70]
  assign _T_397 = _T_396[1]; // @[Shift.scala 12:21]
  assign _T_398 = _T_395[7:0]; // @[Shift.scala 64:52]
  assign _T_400 = {_T_398,2'h0}; // @[Cat.scala 29:58]
  assign _T_401 = _T_397 ? _T_400 : _T_395; // @[Shift.scala 64:27]
  assign _T_402 = _T_396[0:0]; // @[Shift.scala 66:70]
  assign _T_404 = _T_401[8:0]; // @[Shift.scala 64:52]
  assign _T_405 = {_T_404,1'h0}; // @[Cat.scala 29:58]
  assign _T_406 = _T_402 ? _T_405 : _T_401; // @[Shift.scala 64:27]
  assign _T_407 = _T_383 ? _T_406 : 10'h0; // @[Shift.scala 16:10]
  assign _T_408 = _T_407[9:9]; // @[convert.scala 23:34]
  assign decC_fraction = _T_407[8:0]; // @[convert.scala 24:34]
  assign _T_410 = _T_295 == 1'h0; // @[convert.scala 25:26]
  assign _T_412 = _T_295 ? _T_381 : _T_380; // @[convert.scala 25:42]
  assign _T_415 = ~ _T_408; // @[convert.scala 26:67]
  assign _T_416 = _T_293 ? _T_415 : _T_408; // @[convert.scala 26:51]
  assign _T_417 = {_T_410,_T_412,_T_416}; // @[Cat.scala 29:58]
  assign _T_419 = realC[11:0]; // @[convert.scala 29:56]
  assign _T_420 = _T_419 != 12'h0; // @[convert.scala 29:60]
  assign _T_421 = ~ _T_420; // @[convert.scala 29:41]
  assign decC_isNaR = _T_293 & _T_421; // @[convert.scala 29:39]
  assign _T_424 = _T_293 == 1'h0; // @[convert.scala 30:19]
  assign decC_isZero = _T_424 & _T_421; // @[convert.scala 30:41]
  assign decC_scale = $signed(_T_417); // @[convert.scala 32:24]
  assign _T_432 = decA_isNaR | decB_isNaR; // @[PositFMA.scala 58:30]
  assign outIsNaR = _T_432 | decC_isNaR; // @[PositFMA.scala 58:44]
  assign _T_433 = ~ _T_13; // @[PositFMA.scala 59:34]
  assign _T_434 = ~ decA_isZero; // @[PositFMA.scala 59:47]
  assign _T_435 = _T_433 & _T_434; // @[PositFMA.scala 59:45]
  assign _T_437 = {_T_13,_T_435,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_437); // @[PositFMA.scala 59:76]
  assign _T_438 = ~ _T_153; // @[PositFMA.scala 60:34]
  assign _T_439 = ~ decB_isZero; // @[PositFMA.scala 60:47]
  assign _T_440 = _T_438 & _T_439; // @[PositFMA.scala 60:45]
  assign _T_442 = {_T_153,_T_440,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_442); // @[PositFMA.scala 60:76]
  assign _T_443 = $signed(sigA) * $signed(sigB); // @[PositFMA.scala 61:25]
  assign sigP = $unsigned(_T_443); // @[PositFMA.scala 61:33]
  assign _T_444 = sigP[18:0]; // @[PositFMA.scala 62:29]
  assign _T_445 = _T_444 != 19'h0; // @[PositFMA.scala 62:33]
  assign eqTwo = ~ _T_445; // @[PositFMA.scala 62:19]
  assign _T_446 = sigP[20]; // @[PositFMA.scala 64:29]
  assign _T_447 = sigP[19]; // @[PositFMA.scala 64:56]
  assign _T_448 = ~ _T_447; // @[PositFMA.scala 64:51]
  assign _T_449 = _T_446 & _T_448; // @[PositFMA.scala 64:49]
  assign eqFour = _T_449 & eqTwo; // @[PositFMA.scala 64:76]
  assign _T_450 = sigP[21]; // @[PositFMA.scala 66:23]
  assign geTwo = _T_450 ^ _T_447; // @[PositFMA.scala 66:43]
  assign _T_452 = {eqFour,geTwo}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_452)}; // @[PositFMA.scala 67:38]
  assign mulSign = sigP[21:21]; // @[PositFMA.scala 68:28]
  assign _T_453 = $signed(decA_scale) + $signed(decB_scale); // @[PositFMA.scala 70:30]
  assign _GEN_12 = {{4{expBias[2]}},expBias}; // @[PositFMA.scala 70:44]
  assign _T_455 = $signed(_T_453) + $signed(_GEN_12); // @[PositFMA.scala 70:44]
  assign mulScale = $signed(_T_455); // @[PositFMA.scala 70:44]
  assign _T_456 = sigP[19:0]; // @[PositFMA.scala 73:29]
  assign _T_457 = sigP[18:0]; // @[PositFMA.scala 74:29]
  assign _T_458 = {_T_457, 1'h0}; // @[PositFMA.scala 74:48]
  assign mulSigTmp = geTwo ? _T_456 : _T_458; // @[PositFMA.scala 71:22]
  assign _T_460 = mulSigTmp[19:19]; // @[PositFMA.scala 78:39]
  assign _T_461 = _T_460 | eqFour; // @[PositFMA.scala 78:43]
  assign _T_462 = mulSigTmp[18:0]; // @[PositFMA.scala 79:39]
  assign mulSig = {mulSign,_T_461,_T_462}; // @[Cat.scala 29:58]
  assign _T_488 = ~ addSign_phase2; // @[PositFMA.scala 108:29]
  assign _T_489 = ~ addZero_phase2; // @[PositFMA.scala 108:47]
  assign _T_490 = _T_488 & _T_489; // @[PositFMA.scala 108:45]
  assign extAddSig = {addSign_phase2,_T_490,addFrac_phase2,10'h0}; // @[Cat.scala 29:58]
  assign _GEN_13 = {{1{addScale_phase2[5]}},addScale_phase2}; // @[PositFMA.scala 112:39]
  assign mulGreater = $signed(mulScale_phase2) > $signed(_GEN_13); // @[PositFMA.scala 112:39]
  assign greaterScale = mulGreater ? $signed(mulScale_phase2) : $signed({{1{addScale_phase2[5]}},addScale_phase2}); // @[PositFMA.scala 113:26]
  assign smallerScale = mulGreater ? $signed({{1{addScale_phase2[5]}},addScale_phase2}) : $signed(mulScale_phase2); // @[PositFMA.scala 114:26]
  assign _T_494 = $signed(greaterScale) - $signed(smallerScale); // @[PositFMA.scala 115:36]
  assign scaleDiff = $signed(_T_494); // @[PositFMA.scala 115:36]
  assign greaterSig = mulGreater ? mulSig_phase2 : extAddSig; // @[PositFMA.scala 116:26]
  assign smallerSigTmp = mulGreater ? extAddSig : mulSig_phase2; // @[PositFMA.scala 117:26]
  assign _T_495 = $unsigned(scaleDiff); // @[PositFMA.scala 118:69]
  assign _T_496 = _T_495 < 7'h15; // @[Shift.scala 39:24]
  assign _T_497 = _T_495[4:0]; // @[Shift.scala 40:44]
  assign _T_498 = smallerSigTmp[20:16]; // @[Shift.scala 90:30]
  assign _T_499 = smallerSigTmp[15:0]; // @[Shift.scala 90:48]
  assign _T_500 = _T_499 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_14 = {{4'd0}, _T_500}; // @[Shift.scala 90:39]
  assign _T_501 = _T_498 | _GEN_14; // @[Shift.scala 90:39]
  assign _T_502 = _T_497[4]; // @[Shift.scala 12:21]
  assign _T_503 = smallerSigTmp[20]; // @[Shift.scala 12:21]
  assign _T_505 = _T_503 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_506 = {_T_505,_T_501}; // @[Cat.scala 29:58]
  assign _T_507 = _T_502 ? _T_506 : smallerSigTmp; // @[Shift.scala 91:22]
  assign _T_508 = _T_497[3:0]; // @[Shift.scala 92:77]
  assign _T_509 = _T_507[20:8]; // @[Shift.scala 90:30]
  assign _T_510 = _T_507[7:0]; // @[Shift.scala 90:48]
  assign _T_511 = _T_510 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_15 = {{12'd0}, _T_511}; // @[Shift.scala 90:39]
  assign _T_512 = _T_509 | _GEN_15; // @[Shift.scala 90:39]
  assign _T_513 = _T_508[3]; // @[Shift.scala 12:21]
  assign _T_514 = _T_507[20]; // @[Shift.scala 12:21]
  assign _T_516 = _T_514 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_517 = {_T_516,_T_512}; // @[Cat.scala 29:58]
  assign _T_518 = _T_513 ? _T_517 : _T_507; // @[Shift.scala 91:22]
  assign _T_519 = _T_508[2:0]; // @[Shift.scala 92:77]
  assign _T_520 = _T_518[20:4]; // @[Shift.scala 90:30]
  assign _T_521 = _T_518[3:0]; // @[Shift.scala 90:48]
  assign _T_522 = _T_521 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_16 = {{16'd0}, _T_522}; // @[Shift.scala 90:39]
  assign _T_523 = _T_520 | _GEN_16; // @[Shift.scala 90:39]
  assign _T_524 = _T_519[2]; // @[Shift.scala 12:21]
  assign _T_525 = _T_518[20]; // @[Shift.scala 12:21]
  assign _T_527 = _T_525 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_528 = {_T_527,_T_523}; // @[Cat.scala 29:58]
  assign _T_529 = _T_524 ? _T_528 : _T_518; // @[Shift.scala 91:22]
  assign _T_530 = _T_519[1:0]; // @[Shift.scala 92:77]
  assign _T_531 = _T_529[20:2]; // @[Shift.scala 90:30]
  assign _T_532 = _T_529[1:0]; // @[Shift.scala 90:48]
  assign _T_533 = _T_532 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_17 = {{18'd0}, _T_533}; // @[Shift.scala 90:39]
  assign _T_534 = _T_531 | _GEN_17; // @[Shift.scala 90:39]
  assign _T_535 = _T_530[1]; // @[Shift.scala 12:21]
  assign _T_536 = _T_529[20]; // @[Shift.scala 12:21]
  assign _T_538 = _T_536 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_539 = {_T_538,_T_534}; // @[Cat.scala 29:58]
  assign _T_540 = _T_535 ? _T_539 : _T_529; // @[Shift.scala 91:22]
  assign _T_541 = _T_530[0:0]; // @[Shift.scala 92:77]
  assign _T_542 = _T_540[20:1]; // @[Shift.scala 90:30]
  assign _T_543 = _T_540[0:0]; // @[Shift.scala 90:48]
  assign _GEN_18 = {{19'd0}, _T_543}; // @[Shift.scala 90:39]
  assign _T_545 = _T_542 | _GEN_18; // @[Shift.scala 90:39]
  assign _T_547 = _T_540[20]; // @[Shift.scala 12:21]
  assign _T_548 = {_T_547,_T_545}; // @[Cat.scala 29:58]
  assign _T_549 = _T_541 ? _T_548 : _T_540; // @[Shift.scala 91:22]
  assign _T_552 = _T_503 ? 21'h1fffff : 21'h0; // @[Bitwise.scala 71:12]
  assign smallerSig = _T_496 ? _T_549 : _T_552; // @[Shift.scala 39:10]
  assign rawSumSig = greaterSig + smallerSig; // @[PositFMA.scala 119:34]
  assign _T_553 = mulSig_phase2[20:20]; // @[PositFMA.scala 120:42]
  assign _T_554 = _T_553 ^ addSign_phase2; // @[PositFMA.scala 120:46]
  assign _T_555 = rawSumSig[21:21]; // @[PositFMA.scala 120:79]
  assign sumSign = _T_554 ^ _T_555; // @[PositFMA.scala 120:63]
  assign _T_557 = greaterSig + smallerSig; // @[PositFMA.scala 121:50]
  assign signSumSig = {sumSign,_T_557}; // @[Cat.scala 29:58]
  assign _T_558 = signSumSig[21:1]; // @[PositFMA.scala 125:33]
  assign _T_559 = signSumSig[20:0]; // @[PositFMA.scala 125:68]
  assign sumXor = _T_558 ^ _T_559; // @[PositFMA.scala 125:51]
  assign _T_560 = sumXor[20:5]; // @[LZD.scala 43:32]
  assign _T_561 = _T_560[15:8]; // @[LZD.scala 43:32]
  assign _T_562 = _T_561[7:4]; // @[LZD.scala 43:32]
  assign _T_563 = _T_562[3:2]; // @[LZD.scala 43:32]
  assign _T_564 = _T_563 != 2'h0; // @[LZD.scala 39:14]
  assign _T_565 = _T_563[1]; // @[LZD.scala 39:21]
  assign _T_566 = _T_563[0]; // @[LZD.scala 39:30]
  assign _T_567 = ~ _T_566; // @[LZD.scala 39:27]
  assign _T_568 = _T_565 | _T_567; // @[LZD.scala 39:25]
  assign _T_569 = {_T_564,_T_568}; // @[Cat.scala 29:58]
  assign _T_570 = _T_562[1:0]; // @[LZD.scala 44:32]
  assign _T_571 = _T_570 != 2'h0; // @[LZD.scala 39:14]
  assign _T_572 = _T_570[1]; // @[LZD.scala 39:21]
  assign _T_573 = _T_570[0]; // @[LZD.scala 39:30]
  assign _T_574 = ~ _T_573; // @[LZD.scala 39:27]
  assign _T_575 = _T_572 | _T_574; // @[LZD.scala 39:25]
  assign _T_576 = {_T_571,_T_575}; // @[Cat.scala 29:58]
  assign _T_577 = _T_569[1]; // @[Shift.scala 12:21]
  assign _T_578 = _T_576[1]; // @[Shift.scala 12:21]
  assign _T_579 = _T_577 | _T_578; // @[LZD.scala 49:16]
  assign _T_580 = ~ _T_578; // @[LZD.scala 49:27]
  assign _T_581 = _T_577 | _T_580; // @[LZD.scala 49:25]
  assign _T_582 = _T_569[0:0]; // @[LZD.scala 49:47]
  assign _T_583 = _T_576[0:0]; // @[LZD.scala 49:59]
  assign _T_584 = _T_577 ? _T_582 : _T_583; // @[LZD.scala 49:35]
  assign _T_586 = {_T_579,_T_581,_T_584}; // @[Cat.scala 29:58]
  assign _T_587 = _T_561[3:0]; // @[LZD.scala 44:32]
  assign _T_588 = _T_587[3:2]; // @[LZD.scala 43:32]
  assign _T_589 = _T_588 != 2'h0; // @[LZD.scala 39:14]
  assign _T_590 = _T_588[1]; // @[LZD.scala 39:21]
  assign _T_591 = _T_588[0]; // @[LZD.scala 39:30]
  assign _T_592 = ~ _T_591; // @[LZD.scala 39:27]
  assign _T_593 = _T_590 | _T_592; // @[LZD.scala 39:25]
  assign _T_594 = {_T_589,_T_593}; // @[Cat.scala 29:58]
  assign _T_595 = _T_587[1:0]; // @[LZD.scala 44:32]
  assign _T_596 = _T_595 != 2'h0; // @[LZD.scala 39:14]
  assign _T_597 = _T_595[1]; // @[LZD.scala 39:21]
  assign _T_598 = _T_595[0]; // @[LZD.scala 39:30]
  assign _T_599 = ~ _T_598; // @[LZD.scala 39:27]
  assign _T_600 = _T_597 | _T_599; // @[LZD.scala 39:25]
  assign _T_601 = {_T_596,_T_600}; // @[Cat.scala 29:58]
  assign _T_602 = _T_594[1]; // @[Shift.scala 12:21]
  assign _T_603 = _T_601[1]; // @[Shift.scala 12:21]
  assign _T_604 = _T_602 | _T_603; // @[LZD.scala 49:16]
  assign _T_605 = ~ _T_603; // @[LZD.scala 49:27]
  assign _T_606 = _T_602 | _T_605; // @[LZD.scala 49:25]
  assign _T_607 = _T_594[0:0]; // @[LZD.scala 49:47]
  assign _T_608 = _T_601[0:0]; // @[LZD.scala 49:59]
  assign _T_609 = _T_602 ? _T_607 : _T_608; // @[LZD.scala 49:35]
  assign _T_611 = {_T_604,_T_606,_T_609}; // @[Cat.scala 29:58]
  assign _T_612 = _T_586[2]; // @[Shift.scala 12:21]
  assign _T_613 = _T_611[2]; // @[Shift.scala 12:21]
  assign _T_614 = _T_612 | _T_613; // @[LZD.scala 49:16]
  assign _T_615 = ~ _T_613; // @[LZD.scala 49:27]
  assign _T_616 = _T_612 | _T_615; // @[LZD.scala 49:25]
  assign _T_617 = _T_586[1:0]; // @[LZD.scala 49:47]
  assign _T_618 = _T_611[1:0]; // @[LZD.scala 49:59]
  assign _T_619 = _T_612 ? _T_617 : _T_618; // @[LZD.scala 49:35]
  assign _T_621 = {_T_614,_T_616,_T_619}; // @[Cat.scala 29:58]
  assign _T_622 = _T_560[7:0]; // @[LZD.scala 44:32]
  assign _T_623 = _T_622[7:4]; // @[LZD.scala 43:32]
  assign _T_624 = _T_623[3:2]; // @[LZD.scala 43:32]
  assign _T_625 = _T_624 != 2'h0; // @[LZD.scala 39:14]
  assign _T_626 = _T_624[1]; // @[LZD.scala 39:21]
  assign _T_627 = _T_624[0]; // @[LZD.scala 39:30]
  assign _T_628 = ~ _T_627; // @[LZD.scala 39:27]
  assign _T_629 = _T_626 | _T_628; // @[LZD.scala 39:25]
  assign _T_630 = {_T_625,_T_629}; // @[Cat.scala 29:58]
  assign _T_631 = _T_623[1:0]; // @[LZD.scala 44:32]
  assign _T_632 = _T_631 != 2'h0; // @[LZD.scala 39:14]
  assign _T_633 = _T_631[1]; // @[LZD.scala 39:21]
  assign _T_634 = _T_631[0]; // @[LZD.scala 39:30]
  assign _T_635 = ~ _T_634; // @[LZD.scala 39:27]
  assign _T_636 = _T_633 | _T_635; // @[LZD.scala 39:25]
  assign _T_637 = {_T_632,_T_636}; // @[Cat.scala 29:58]
  assign _T_638 = _T_630[1]; // @[Shift.scala 12:21]
  assign _T_639 = _T_637[1]; // @[Shift.scala 12:21]
  assign _T_640 = _T_638 | _T_639; // @[LZD.scala 49:16]
  assign _T_641 = ~ _T_639; // @[LZD.scala 49:27]
  assign _T_642 = _T_638 | _T_641; // @[LZD.scala 49:25]
  assign _T_643 = _T_630[0:0]; // @[LZD.scala 49:47]
  assign _T_644 = _T_637[0:0]; // @[LZD.scala 49:59]
  assign _T_645 = _T_638 ? _T_643 : _T_644; // @[LZD.scala 49:35]
  assign _T_647 = {_T_640,_T_642,_T_645}; // @[Cat.scala 29:58]
  assign _T_648 = _T_622[3:0]; // @[LZD.scala 44:32]
  assign _T_649 = _T_648[3:2]; // @[LZD.scala 43:32]
  assign _T_650 = _T_649 != 2'h0; // @[LZD.scala 39:14]
  assign _T_651 = _T_649[1]; // @[LZD.scala 39:21]
  assign _T_652 = _T_649[0]; // @[LZD.scala 39:30]
  assign _T_653 = ~ _T_652; // @[LZD.scala 39:27]
  assign _T_654 = _T_651 | _T_653; // @[LZD.scala 39:25]
  assign _T_655 = {_T_650,_T_654}; // @[Cat.scala 29:58]
  assign _T_656 = _T_648[1:0]; // @[LZD.scala 44:32]
  assign _T_657 = _T_656 != 2'h0; // @[LZD.scala 39:14]
  assign _T_658 = _T_656[1]; // @[LZD.scala 39:21]
  assign _T_659 = _T_656[0]; // @[LZD.scala 39:30]
  assign _T_660 = ~ _T_659; // @[LZD.scala 39:27]
  assign _T_661 = _T_658 | _T_660; // @[LZD.scala 39:25]
  assign _T_662 = {_T_657,_T_661}; // @[Cat.scala 29:58]
  assign _T_663 = _T_655[1]; // @[Shift.scala 12:21]
  assign _T_664 = _T_662[1]; // @[Shift.scala 12:21]
  assign _T_665 = _T_663 | _T_664; // @[LZD.scala 49:16]
  assign _T_666 = ~ _T_664; // @[LZD.scala 49:27]
  assign _T_667 = _T_663 | _T_666; // @[LZD.scala 49:25]
  assign _T_668 = _T_655[0:0]; // @[LZD.scala 49:47]
  assign _T_669 = _T_662[0:0]; // @[LZD.scala 49:59]
  assign _T_670 = _T_663 ? _T_668 : _T_669; // @[LZD.scala 49:35]
  assign _T_672 = {_T_665,_T_667,_T_670}; // @[Cat.scala 29:58]
  assign _T_673 = _T_647[2]; // @[Shift.scala 12:21]
  assign _T_674 = _T_672[2]; // @[Shift.scala 12:21]
  assign _T_675 = _T_673 | _T_674; // @[LZD.scala 49:16]
  assign _T_676 = ~ _T_674; // @[LZD.scala 49:27]
  assign _T_677 = _T_673 | _T_676; // @[LZD.scala 49:25]
  assign _T_678 = _T_647[1:0]; // @[LZD.scala 49:47]
  assign _T_679 = _T_672[1:0]; // @[LZD.scala 49:59]
  assign _T_680 = _T_673 ? _T_678 : _T_679; // @[LZD.scala 49:35]
  assign _T_682 = {_T_675,_T_677,_T_680}; // @[Cat.scala 29:58]
  assign _T_683 = _T_621[3]; // @[Shift.scala 12:21]
  assign _T_684 = _T_682[3]; // @[Shift.scala 12:21]
  assign _T_685 = _T_683 | _T_684; // @[LZD.scala 49:16]
  assign _T_686 = ~ _T_684; // @[LZD.scala 49:27]
  assign _T_687 = _T_683 | _T_686; // @[LZD.scala 49:25]
  assign _T_688 = _T_621[2:0]; // @[LZD.scala 49:47]
  assign _T_689 = _T_682[2:0]; // @[LZD.scala 49:59]
  assign _T_690 = _T_683 ? _T_688 : _T_689; // @[LZD.scala 49:35]
  assign _T_692 = {_T_685,_T_687,_T_690}; // @[Cat.scala 29:58]
  assign _T_693 = sumXor[4:0]; // @[LZD.scala 44:32]
  assign _T_694 = _T_693[4:1]; // @[LZD.scala 43:32]
  assign _T_695 = _T_694[3:2]; // @[LZD.scala 43:32]
  assign _T_696 = _T_695 != 2'h0; // @[LZD.scala 39:14]
  assign _T_697 = _T_695[1]; // @[LZD.scala 39:21]
  assign _T_698 = _T_695[0]; // @[LZD.scala 39:30]
  assign _T_699 = ~ _T_698; // @[LZD.scala 39:27]
  assign _T_700 = _T_697 | _T_699; // @[LZD.scala 39:25]
  assign _T_701 = {_T_696,_T_700}; // @[Cat.scala 29:58]
  assign _T_702 = _T_694[1:0]; // @[LZD.scala 44:32]
  assign _T_703 = _T_702 != 2'h0; // @[LZD.scala 39:14]
  assign _T_704 = _T_702[1]; // @[LZD.scala 39:21]
  assign _T_705 = _T_702[0]; // @[LZD.scala 39:30]
  assign _T_706 = ~ _T_705; // @[LZD.scala 39:27]
  assign _T_707 = _T_704 | _T_706; // @[LZD.scala 39:25]
  assign _T_708 = {_T_703,_T_707}; // @[Cat.scala 29:58]
  assign _T_709 = _T_701[1]; // @[Shift.scala 12:21]
  assign _T_710 = _T_708[1]; // @[Shift.scala 12:21]
  assign _T_711 = _T_709 | _T_710; // @[LZD.scala 49:16]
  assign _T_712 = ~ _T_710; // @[LZD.scala 49:27]
  assign _T_713 = _T_709 | _T_712; // @[LZD.scala 49:25]
  assign _T_714 = _T_701[0:0]; // @[LZD.scala 49:47]
  assign _T_715 = _T_708[0:0]; // @[LZD.scala 49:59]
  assign _T_716 = _T_709 ? _T_714 : _T_715; // @[LZD.scala 49:35]
  assign _T_718 = {_T_711,_T_713,_T_716}; // @[Cat.scala 29:58]
  assign _T_719 = _T_693[0:0]; // @[LZD.scala 44:32]
  assign _T_721 = _T_718[2]; // @[Shift.scala 12:21]
  assign _T_723 = {1'h1,_T_719}; // @[Cat.scala 29:58]
  assign _T_724 = _T_718[1:0]; // @[LZD.scala 55:32]
  assign _T_725 = _T_721 ? _T_724 : _T_723; // @[LZD.scala 55:20]
  assign _T_727 = _T_692[4]; // @[Shift.scala 12:21]
  assign _T_729 = {1'h1,_T_721,_T_725}; // @[Cat.scala 29:58]
  assign _T_730 = _T_692[3:0]; // @[LZD.scala 55:32]
  assign _T_731 = _T_727 ? _T_730 : _T_729; // @[LZD.scala 55:20]
  assign sumLZD = {_T_727,_T_731}; // @[Cat.scala 29:58]
  assign shiftValue = ~ sumLZD; // @[PositFMA.scala 127:24]
  assign _T_732 = signSumSig[19:0]; // @[PositFMA.scala 128:38]
  assign _T_733 = shiftValue < 5'h14; // @[Shift.scala 16:24]
  assign _T_735 = shiftValue[4]; // @[Shift.scala 12:21]
  assign _T_736 = _T_732[3:0]; // @[Shift.scala 64:52]
  assign _T_738 = {_T_736,16'h0}; // @[Cat.scala 29:58]
  assign _T_739 = _T_735 ? _T_738 : _T_732; // @[Shift.scala 64:27]
  assign _T_740 = shiftValue[3:0]; // @[Shift.scala 66:70]
  assign _T_741 = _T_740[3]; // @[Shift.scala 12:21]
  assign _T_742 = _T_739[11:0]; // @[Shift.scala 64:52]
  assign _T_744 = {_T_742,8'h0}; // @[Cat.scala 29:58]
  assign _T_745 = _T_741 ? _T_744 : _T_739; // @[Shift.scala 64:27]
  assign _T_746 = _T_740[2:0]; // @[Shift.scala 66:70]
  assign _T_747 = _T_746[2]; // @[Shift.scala 12:21]
  assign _T_748 = _T_745[15:0]; // @[Shift.scala 64:52]
  assign _T_750 = {_T_748,4'h0}; // @[Cat.scala 29:58]
  assign _T_751 = _T_747 ? _T_750 : _T_745; // @[Shift.scala 64:27]
  assign _T_752 = _T_746[1:0]; // @[Shift.scala 66:70]
  assign _T_753 = _T_752[1]; // @[Shift.scala 12:21]
  assign _T_754 = _T_751[17:0]; // @[Shift.scala 64:52]
  assign _T_756 = {_T_754,2'h0}; // @[Cat.scala 29:58]
  assign _T_757 = _T_753 ? _T_756 : _T_751; // @[Shift.scala 64:27]
  assign _T_758 = _T_752[0:0]; // @[Shift.scala 66:70]
  assign _T_760 = _T_757[18:0]; // @[Shift.scala 64:52]
  assign _T_761 = {_T_760,1'h0}; // @[Cat.scala 29:58]
  assign _T_762 = _T_758 ? _T_761 : _T_757; // @[Shift.scala 64:27]
  assign normalFracTmp = _T_733 ? _T_762 : 20'h0; // @[Shift.scala 16:10]
  assign _T_764 = $signed(greaterScale) + $signed(7'sh2); // @[PositFMA.scala 131:36]
  assign _T_765 = $signed(_T_764); // @[PositFMA.scala 131:36]
  assign _T_766 = {1'h1,_T_727,_T_731}; // @[Cat.scala 29:58]
  assign _T_767 = $signed(_T_766); // @[PositFMA.scala 131:61]
  assign _GEN_19 = {{1{_T_767[5]}},_T_767}; // @[PositFMA.scala 131:42]
  assign _T_769 = $signed(_T_765) + $signed(_GEN_19); // @[PositFMA.scala 131:42]
  assign sumScale = $signed(_T_769); // @[PositFMA.scala 131:42]
  assign sumFrac = normalFracTmp[19:11]; // @[PositFMA.scala 132:41]
  assign grsTmp = normalFracTmp[10:0]; // @[PositFMA.scala 135:41]
  assign _T_770 = grsTmp[10:9]; // @[PositFMA.scala 138:40]
  assign _T_771 = grsTmp[8:0]; // @[PositFMA.scala 138:56]
  assign _T_772 = _T_771 != 9'h0; // @[PositFMA.scala 138:60]
  assign underflow = $signed(sumScale) < $signed(-7'sh16); // @[PositFMA.scala 145:32]
  assign overflow = $signed(sumScale) > $signed(7'sh16); // @[PositFMA.scala 146:32]
  assign _T_773 = signSumSig != 22'h0; // @[PositFMA.scala 155:32]
  assign decF_isZero = ~ _T_773; // @[PositFMA.scala 155:20]
  assign _T_775 = underflow ? $signed(-7'sh16) : $signed(sumScale); // @[Mux.scala 87:16]
  assign _T_776 = overflow ? $signed(7'sh16) : $signed(_T_775); // @[Mux.scala 87:16]
  assign _GEN_20 = _T_776[5:0]; // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  assign decF_scale = $signed(_GEN_20); // @[PositFMA.scala 152:18 PositFMA.scala 158:17]
  assign _T_777 = decF_scale[0]; // @[convert.scala 46:61]
  assign _T_778 = ~ _T_777; // @[convert.scala 46:52]
  assign _T_780 = sumSign ? _T_778 : _T_777; // @[convert.scala 46:42]
  assign _T_781 = decF_scale[5:1]; // @[convert.scala 48:34]
  assign _T_782 = _T_781[4:4]; // @[convert.scala 49:36]
  assign _T_784 = ~ _T_781; // @[convert.scala 50:36]
  assign _T_785 = $signed(_T_784); // @[convert.scala 50:36]
  assign _T_786 = _T_782 ? $signed(_T_785) : $signed(_T_781); // @[convert.scala 50:28]
  assign _T_787 = _T_782 ^ sumSign; // @[convert.scala 51:31]
  assign _T_788 = ~ _T_787; // @[convert.scala 52:43]
  assign _T_792 = {_T_788,_T_787,_T_780,sumFrac,_T_770,_T_772}; // @[Cat.scala 29:58]
  assign _T_793 = $unsigned(_T_786); // @[Shift.scala 39:17]
  assign _T_794 = _T_793 < 5'hf; // @[Shift.scala 39:24]
  assign _T_795 = _T_786[3:0]; // @[Shift.scala 40:44]
  assign _T_796 = _T_792[14:8]; // @[Shift.scala 90:30]
  assign _T_797 = _T_792[7:0]; // @[Shift.scala 90:48]
  assign _T_798 = _T_797 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{6'd0}, _T_798}; // @[Shift.scala 90:39]
  assign _T_799 = _T_796 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_800 = _T_795[3]; // @[Shift.scala 12:21]
  assign _T_801 = _T_792[14]; // @[Shift.scala 12:21]
  assign _T_803 = _T_801 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_804 = {_T_803,_T_799}; // @[Cat.scala 29:58]
  assign _T_805 = _T_800 ? _T_804 : _T_792; // @[Shift.scala 91:22]
  assign _T_806 = _T_795[2:0]; // @[Shift.scala 92:77]
  assign _T_807 = _T_805[14:4]; // @[Shift.scala 90:30]
  assign _T_808 = _T_805[3:0]; // @[Shift.scala 90:48]
  assign _T_809 = _T_808 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{10'd0}, _T_809}; // @[Shift.scala 90:39]
  assign _T_810 = _T_807 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_811 = _T_806[2]; // @[Shift.scala 12:21]
  assign _T_812 = _T_805[14]; // @[Shift.scala 12:21]
  assign _T_814 = _T_812 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_815 = {_T_814,_T_810}; // @[Cat.scala 29:58]
  assign _T_816 = _T_811 ? _T_815 : _T_805; // @[Shift.scala 91:22]
  assign _T_817 = _T_806[1:0]; // @[Shift.scala 92:77]
  assign _T_818 = _T_816[14:2]; // @[Shift.scala 90:30]
  assign _T_819 = _T_816[1:0]; // @[Shift.scala 90:48]
  assign _T_820 = _T_819 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_23 = {{12'd0}, _T_820}; // @[Shift.scala 90:39]
  assign _T_821 = _T_818 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_822 = _T_817[1]; // @[Shift.scala 12:21]
  assign _T_823 = _T_816[14]; // @[Shift.scala 12:21]
  assign _T_825 = _T_823 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_826 = {_T_825,_T_821}; // @[Cat.scala 29:58]
  assign _T_827 = _T_822 ? _T_826 : _T_816; // @[Shift.scala 91:22]
  assign _T_828 = _T_817[0:0]; // @[Shift.scala 92:77]
  assign _T_829 = _T_827[14:1]; // @[Shift.scala 90:30]
  assign _T_830 = _T_827[0:0]; // @[Shift.scala 90:48]
  assign _GEN_24 = {{13'd0}, _T_830}; // @[Shift.scala 90:39]
  assign _T_832 = _T_829 | _GEN_24; // @[Shift.scala 90:39]
  assign _T_834 = _T_827[14]; // @[Shift.scala 12:21]
  assign _T_835 = {_T_834,_T_832}; // @[Cat.scala 29:58]
  assign _T_836 = _T_828 ? _T_835 : _T_827; // @[Shift.scala 91:22]
  assign _T_839 = _T_801 ? 15'h7fff : 15'h0; // @[Bitwise.scala 71:12]
  assign _T_840 = _T_794 ? _T_836 : _T_839; // @[Shift.scala 39:10]
  assign _T_841 = _T_840[3]; // @[convert.scala 55:31]
  assign _T_842 = _T_840[2]; // @[convert.scala 56:31]
  assign _T_843 = _T_840[1]; // @[convert.scala 57:31]
  assign _T_844 = _T_840[0]; // @[convert.scala 58:31]
  assign _T_845 = _T_840[14:3]; // @[convert.scala 59:69]
  assign _T_846 = _T_845 != 12'h0; // @[convert.scala 59:81]
  assign _T_847 = ~ _T_846; // @[convert.scala 59:50]
  assign _T_849 = _T_845 == 12'hfff; // @[convert.scala 60:81]
  assign _T_850 = _T_841 | _T_843; // @[convert.scala 61:44]
  assign _T_851 = _T_850 | _T_844; // @[convert.scala 61:52]
  assign _T_852 = _T_842 & _T_851; // @[convert.scala 61:36]
  assign _T_853 = ~ _T_849; // @[convert.scala 62:63]
  assign _T_854 = _T_853 & _T_852; // @[convert.scala 62:103]
  assign _T_855 = _T_847 | _T_854; // @[convert.scala 62:60]
  assign _GEN_25 = {{11'd0}, _T_855}; // @[convert.scala 63:56]
  assign _T_858 = _T_845 + _GEN_25; // @[convert.scala 63:56]
  assign _T_859 = {sumSign,_T_858}; // @[Cat.scala 29:58]
  assign io_F = _T_867; // @[PositFMA.scala 175:15]
  assign io_outValid = _T_863; // @[PositFMA.scala 174:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  outIsNaR_phase2 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mulSig_phase2 = _RAND_1[20:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  addFrac_phase2 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mulScale_phase2 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addScale_phase2 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addSign_phase2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addZero_phase2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inValid_phase2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_863 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_867 = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_inValid) begin
      outIsNaR_phase2 <= outIsNaR;
    end
    if (io_inValid) begin
      mulSig_phase2 <= mulSig;
    end
    if (io_inValid) begin
      addFrac_phase2 <= decC_fraction;
    end
    if (io_inValid) begin
      mulScale_phase2 <= mulScale;
    end
    if (io_inValid) begin
      addScale_phase2 <= decC_scale;
    end
    if (io_inValid) begin
      addSign_phase2 <= _T_293;
    end
    if (io_inValid) begin
      addZero_phase2 <= decC_isZero;
    end
    if (reset) begin
      inValid_phase2 <= 1'h0;
    end else begin
      inValid_phase2 <= io_inValid;
    end
    if (reset) begin
      _T_863 <= 1'h0;
    end else begin
      _T_863 <= inValid_phase2;
    end
    if (inValid_phase2) begin
      if (outIsNaR_phase2) begin
        _T_867 <= 13'h1000;
      end else begin
        if (decF_isZero) begin
          _T_867 <= 13'h0;
        end else begin
          _T_867 <= _T_859;
        end
      end
    end
  end
endmodule
