module QuireToPosit30_8_2(
  input          clock,
  input          reset,
  input          io_inValid,
  input  [127:0] io_quireIn,
  output [7:0]   io_positOut,
  output         io_outValid
);
  wire [126:0] _T; // @[QuireToPosit.scala 47:43]
  wire  _T_1; // @[QuireToPosit.scala 47:47]
  wire  tailIsZero; // @[QuireToPosit.scala 47:27]
  wire  _T_2; // @[QuireToPosit.scala 49:45]
  wire  outRawFloat_isNaR; // @[QuireToPosit.scala 49:49]
  wire  _T_5; // @[QuireToPosit.scala 50:31]
  wire  outRawFloat_isZero; // @[QuireToPosit.scala 50:51]
  wire [126:0] _T_8; // @[QuireToPosit.scala 58:41]
  wire [126:0] _T_9; // @[QuireToPosit.scala 58:68]
  wire [126:0] quireXOR; // @[QuireToPosit.scala 58:56]
  wire [63:0] _T_10; // @[LZD.scala 43:32]
  wire [31:0] _T_11; // @[LZD.scala 43:32]
  wire [15:0] _T_12; // @[LZD.scala 43:32]
  wire [7:0] _T_13; // @[LZD.scala 43:32]
  wire [3:0] _T_14; // @[LZD.scala 43:32]
  wire [1:0] _T_15; // @[LZD.scala 43:32]
  wire  _T_16; // @[LZD.scala 39:14]
  wire  _T_17; // @[LZD.scala 39:21]
  wire  _T_18; // @[LZD.scala 39:30]
  wire  _T_19; // @[LZD.scala 39:27]
  wire  _T_20; // @[LZD.scala 39:25]
  wire [1:0] _T_21; // @[Cat.scala 29:58]
  wire [1:0] _T_22; // @[LZD.scala 44:32]
  wire  _T_23; // @[LZD.scala 39:14]
  wire  _T_24; // @[LZD.scala 39:21]
  wire  _T_25; // @[LZD.scala 39:30]
  wire  _T_26; // @[LZD.scala 39:27]
  wire  _T_27; // @[LZD.scala 39:25]
  wire [1:0] _T_28; // @[Cat.scala 29:58]
  wire  _T_29; // @[Shift.scala 12:21]
  wire  _T_30; // @[Shift.scala 12:21]
  wire  _T_31; // @[LZD.scala 49:16]
  wire  _T_32; // @[LZD.scala 49:27]
  wire  _T_33; // @[LZD.scala 49:25]
  wire  _T_34; // @[LZD.scala 49:47]
  wire  _T_35; // @[LZD.scala 49:59]
  wire  _T_36; // @[LZD.scala 49:35]
  wire [2:0] _T_38; // @[Cat.scala 29:58]
  wire [3:0] _T_39; // @[LZD.scala 44:32]
  wire [1:0] _T_40; // @[LZD.scala 43:32]
  wire  _T_41; // @[LZD.scala 39:14]
  wire  _T_42; // @[LZD.scala 39:21]
  wire  _T_43; // @[LZD.scala 39:30]
  wire  _T_44; // @[LZD.scala 39:27]
  wire  _T_45; // @[LZD.scala 39:25]
  wire [1:0] _T_46; // @[Cat.scala 29:58]
  wire [1:0] _T_47; // @[LZD.scala 44:32]
  wire  _T_48; // @[LZD.scala 39:14]
  wire  _T_49; // @[LZD.scala 39:21]
  wire  _T_50; // @[LZD.scala 39:30]
  wire  _T_51; // @[LZD.scala 39:27]
  wire  _T_52; // @[LZD.scala 39:25]
  wire [1:0] _T_53; // @[Cat.scala 29:58]
  wire  _T_54; // @[Shift.scala 12:21]
  wire  _T_55; // @[Shift.scala 12:21]
  wire  _T_56; // @[LZD.scala 49:16]
  wire  _T_57; // @[LZD.scala 49:27]
  wire  _T_58; // @[LZD.scala 49:25]
  wire  _T_59; // @[LZD.scala 49:47]
  wire  _T_60; // @[LZD.scala 49:59]
  wire  _T_61; // @[LZD.scala 49:35]
  wire [2:0] _T_63; // @[Cat.scala 29:58]
  wire  _T_64; // @[Shift.scala 12:21]
  wire  _T_65; // @[Shift.scala 12:21]
  wire  _T_66; // @[LZD.scala 49:16]
  wire  _T_67; // @[LZD.scala 49:27]
  wire  _T_68; // @[LZD.scala 49:25]
  wire [1:0] _T_69; // @[LZD.scala 49:47]
  wire [1:0] _T_70; // @[LZD.scala 49:59]
  wire [1:0] _T_71; // @[LZD.scala 49:35]
  wire [3:0] _T_73; // @[Cat.scala 29:58]
  wire [7:0] _T_74; // @[LZD.scala 44:32]
  wire [3:0] _T_75; // @[LZD.scala 43:32]
  wire [1:0] _T_76; // @[LZD.scala 43:32]
  wire  _T_77; // @[LZD.scala 39:14]
  wire  _T_78; // @[LZD.scala 39:21]
  wire  _T_79; // @[LZD.scala 39:30]
  wire  _T_80; // @[LZD.scala 39:27]
  wire  _T_81; // @[LZD.scala 39:25]
  wire [1:0] _T_82; // @[Cat.scala 29:58]
  wire [1:0] _T_83; // @[LZD.scala 44:32]
  wire  _T_84; // @[LZD.scala 39:14]
  wire  _T_85; // @[LZD.scala 39:21]
  wire  _T_86; // @[LZD.scala 39:30]
  wire  _T_87; // @[LZD.scala 39:27]
  wire  _T_88; // @[LZD.scala 39:25]
  wire [1:0] _T_89; // @[Cat.scala 29:58]
  wire  _T_90; // @[Shift.scala 12:21]
  wire  _T_91; // @[Shift.scala 12:21]
  wire  _T_92; // @[LZD.scala 49:16]
  wire  _T_93; // @[LZD.scala 49:27]
  wire  _T_94; // @[LZD.scala 49:25]
  wire  _T_95; // @[LZD.scala 49:47]
  wire  _T_96; // @[LZD.scala 49:59]
  wire  _T_97; // @[LZD.scala 49:35]
  wire [2:0] _T_99; // @[Cat.scala 29:58]
  wire [3:0] _T_100; // @[LZD.scala 44:32]
  wire [1:0] _T_101; // @[LZD.scala 43:32]
  wire  _T_102; // @[LZD.scala 39:14]
  wire  _T_103; // @[LZD.scala 39:21]
  wire  _T_104; // @[LZD.scala 39:30]
  wire  _T_105; // @[LZD.scala 39:27]
  wire  _T_106; // @[LZD.scala 39:25]
  wire [1:0] _T_107; // @[Cat.scala 29:58]
  wire [1:0] _T_108; // @[LZD.scala 44:32]
  wire  _T_109; // @[LZD.scala 39:14]
  wire  _T_110; // @[LZD.scala 39:21]
  wire  _T_111; // @[LZD.scala 39:30]
  wire  _T_112; // @[LZD.scala 39:27]
  wire  _T_113; // @[LZD.scala 39:25]
  wire [1:0] _T_114; // @[Cat.scala 29:58]
  wire  _T_115; // @[Shift.scala 12:21]
  wire  _T_116; // @[Shift.scala 12:21]
  wire  _T_117; // @[LZD.scala 49:16]
  wire  _T_118; // @[LZD.scala 49:27]
  wire  _T_119; // @[LZD.scala 49:25]
  wire  _T_120; // @[LZD.scala 49:47]
  wire  _T_121; // @[LZD.scala 49:59]
  wire  _T_122; // @[LZD.scala 49:35]
  wire [2:0] _T_124; // @[Cat.scala 29:58]
  wire  _T_125; // @[Shift.scala 12:21]
  wire  _T_126; // @[Shift.scala 12:21]
  wire  _T_127; // @[LZD.scala 49:16]
  wire  _T_128; // @[LZD.scala 49:27]
  wire  _T_129; // @[LZD.scala 49:25]
  wire [1:0] _T_130; // @[LZD.scala 49:47]
  wire [1:0] _T_131; // @[LZD.scala 49:59]
  wire [1:0] _T_132; // @[LZD.scala 49:35]
  wire [3:0] _T_134; // @[Cat.scala 29:58]
  wire  _T_135; // @[Shift.scala 12:21]
  wire  _T_136; // @[Shift.scala 12:21]
  wire  _T_137; // @[LZD.scala 49:16]
  wire  _T_138; // @[LZD.scala 49:27]
  wire  _T_139; // @[LZD.scala 49:25]
  wire [2:0] _T_140; // @[LZD.scala 49:47]
  wire [2:0] _T_141; // @[LZD.scala 49:59]
  wire [2:0] _T_142; // @[LZD.scala 49:35]
  wire [4:0] _T_144; // @[Cat.scala 29:58]
  wire [15:0] _T_145; // @[LZD.scala 44:32]
  wire [7:0] _T_146; // @[LZD.scala 43:32]
  wire [3:0] _T_147; // @[LZD.scala 43:32]
  wire [1:0] _T_148; // @[LZD.scala 43:32]
  wire  _T_149; // @[LZD.scala 39:14]
  wire  _T_150; // @[LZD.scala 39:21]
  wire  _T_151; // @[LZD.scala 39:30]
  wire  _T_152; // @[LZD.scala 39:27]
  wire  _T_153; // @[LZD.scala 39:25]
  wire [1:0] _T_154; // @[Cat.scala 29:58]
  wire [1:0] _T_155; // @[LZD.scala 44:32]
  wire  _T_156; // @[LZD.scala 39:14]
  wire  _T_157; // @[LZD.scala 39:21]
  wire  _T_158; // @[LZD.scala 39:30]
  wire  _T_159; // @[LZD.scala 39:27]
  wire  _T_160; // @[LZD.scala 39:25]
  wire [1:0] _T_161; // @[Cat.scala 29:58]
  wire  _T_162; // @[Shift.scala 12:21]
  wire  _T_163; // @[Shift.scala 12:21]
  wire  _T_164; // @[LZD.scala 49:16]
  wire  _T_165; // @[LZD.scala 49:27]
  wire  _T_166; // @[LZD.scala 49:25]
  wire  _T_167; // @[LZD.scala 49:47]
  wire  _T_168; // @[LZD.scala 49:59]
  wire  _T_169; // @[LZD.scala 49:35]
  wire [2:0] _T_171; // @[Cat.scala 29:58]
  wire [3:0] _T_172; // @[LZD.scala 44:32]
  wire [1:0] _T_173; // @[LZD.scala 43:32]
  wire  _T_174; // @[LZD.scala 39:14]
  wire  _T_175; // @[LZD.scala 39:21]
  wire  _T_176; // @[LZD.scala 39:30]
  wire  _T_177; // @[LZD.scala 39:27]
  wire  _T_178; // @[LZD.scala 39:25]
  wire [1:0] _T_179; // @[Cat.scala 29:58]
  wire [1:0] _T_180; // @[LZD.scala 44:32]
  wire  _T_181; // @[LZD.scala 39:14]
  wire  _T_182; // @[LZD.scala 39:21]
  wire  _T_183; // @[LZD.scala 39:30]
  wire  _T_184; // @[LZD.scala 39:27]
  wire  _T_185; // @[LZD.scala 39:25]
  wire [1:0] _T_186; // @[Cat.scala 29:58]
  wire  _T_187; // @[Shift.scala 12:21]
  wire  _T_188; // @[Shift.scala 12:21]
  wire  _T_189; // @[LZD.scala 49:16]
  wire  _T_190; // @[LZD.scala 49:27]
  wire  _T_191; // @[LZD.scala 49:25]
  wire  _T_192; // @[LZD.scala 49:47]
  wire  _T_193; // @[LZD.scala 49:59]
  wire  _T_194; // @[LZD.scala 49:35]
  wire [2:0] _T_196; // @[Cat.scala 29:58]
  wire  _T_197; // @[Shift.scala 12:21]
  wire  _T_198; // @[Shift.scala 12:21]
  wire  _T_199; // @[LZD.scala 49:16]
  wire  _T_200; // @[LZD.scala 49:27]
  wire  _T_201; // @[LZD.scala 49:25]
  wire [1:0] _T_202; // @[LZD.scala 49:47]
  wire [1:0] _T_203; // @[LZD.scala 49:59]
  wire [1:0] _T_204; // @[LZD.scala 49:35]
  wire [3:0] _T_206; // @[Cat.scala 29:58]
  wire [7:0] _T_207; // @[LZD.scala 44:32]
  wire [3:0] _T_208; // @[LZD.scala 43:32]
  wire [1:0] _T_209; // @[LZD.scala 43:32]
  wire  _T_210; // @[LZD.scala 39:14]
  wire  _T_211; // @[LZD.scala 39:21]
  wire  _T_212; // @[LZD.scala 39:30]
  wire  _T_213; // @[LZD.scala 39:27]
  wire  _T_214; // @[LZD.scala 39:25]
  wire [1:0] _T_215; // @[Cat.scala 29:58]
  wire [1:0] _T_216; // @[LZD.scala 44:32]
  wire  _T_217; // @[LZD.scala 39:14]
  wire  _T_218; // @[LZD.scala 39:21]
  wire  _T_219; // @[LZD.scala 39:30]
  wire  _T_220; // @[LZD.scala 39:27]
  wire  _T_221; // @[LZD.scala 39:25]
  wire [1:0] _T_222; // @[Cat.scala 29:58]
  wire  _T_223; // @[Shift.scala 12:21]
  wire  _T_224; // @[Shift.scala 12:21]
  wire  _T_225; // @[LZD.scala 49:16]
  wire  _T_226; // @[LZD.scala 49:27]
  wire  _T_227; // @[LZD.scala 49:25]
  wire  _T_228; // @[LZD.scala 49:47]
  wire  _T_229; // @[LZD.scala 49:59]
  wire  _T_230; // @[LZD.scala 49:35]
  wire [2:0] _T_232; // @[Cat.scala 29:58]
  wire [3:0] _T_233; // @[LZD.scala 44:32]
  wire [1:0] _T_234; // @[LZD.scala 43:32]
  wire  _T_235; // @[LZD.scala 39:14]
  wire  _T_236; // @[LZD.scala 39:21]
  wire  _T_237; // @[LZD.scala 39:30]
  wire  _T_238; // @[LZD.scala 39:27]
  wire  _T_239; // @[LZD.scala 39:25]
  wire [1:0] _T_240; // @[Cat.scala 29:58]
  wire [1:0] _T_241; // @[LZD.scala 44:32]
  wire  _T_242; // @[LZD.scala 39:14]
  wire  _T_243; // @[LZD.scala 39:21]
  wire  _T_244; // @[LZD.scala 39:30]
  wire  _T_245; // @[LZD.scala 39:27]
  wire  _T_246; // @[LZD.scala 39:25]
  wire [1:0] _T_247; // @[Cat.scala 29:58]
  wire  _T_248; // @[Shift.scala 12:21]
  wire  _T_249; // @[Shift.scala 12:21]
  wire  _T_250; // @[LZD.scala 49:16]
  wire  _T_251; // @[LZD.scala 49:27]
  wire  _T_252; // @[LZD.scala 49:25]
  wire  _T_253; // @[LZD.scala 49:47]
  wire  _T_254; // @[LZD.scala 49:59]
  wire  _T_255; // @[LZD.scala 49:35]
  wire [2:0] _T_257; // @[Cat.scala 29:58]
  wire  _T_258; // @[Shift.scala 12:21]
  wire  _T_259; // @[Shift.scala 12:21]
  wire  _T_260; // @[LZD.scala 49:16]
  wire  _T_261; // @[LZD.scala 49:27]
  wire  _T_262; // @[LZD.scala 49:25]
  wire [1:0] _T_263; // @[LZD.scala 49:47]
  wire [1:0] _T_264; // @[LZD.scala 49:59]
  wire [1:0] _T_265; // @[LZD.scala 49:35]
  wire [3:0] _T_267; // @[Cat.scala 29:58]
  wire  _T_268; // @[Shift.scala 12:21]
  wire  _T_269; // @[Shift.scala 12:21]
  wire  _T_270; // @[LZD.scala 49:16]
  wire  _T_271; // @[LZD.scala 49:27]
  wire  _T_272; // @[LZD.scala 49:25]
  wire [2:0] _T_273; // @[LZD.scala 49:47]
  wire [2:0] _T_274; // @[LZD.scala 49:59]
  wire [2:0] _T_275; // @[LZD.scala 49:35]
  wire [4:0] _T_277; // @[Cat.scala 29:58]
  wire  _T_278; // @[Shift.scala 12:21]
  wire  _T_279; // @[Shift.scala 12:21]
  wire  _T_280; // @[LZD.scala 49:16]
  wire  _T_281; // @[LZD.scala 49:27]
  wire  _T_282; // @[LZD.scala 49:25]
  wire [3:0] _T_283; // @[LZD.scala 49:47]
  wire [3:0] _T_284; // @[LZD.scala 49:59]
  wire [3:0] _T_285; // @[LZD.scala 49:35]
  wire [5:0] _T_287; // @[Cat.scala 29:58]
  wire [31:0] _T_288; // @[LZD.scala 44:32]
  wire [15:0] _T_289; // @[LZD.scala 43:32]
  wire [7:0] _T_290; // @[LZD.scala 43:32]
  wire [3:0] _T_291; // @[LZD.scala 43:32]
  wire [1:0] _T_292; // @[LZD.scala 43:32]
  wire  _T_293; // @[LZD.scala 39:14]
  wire  _T_294; // @[LZD.scala 39:21]
  wire  _T_295; // @[LZD.scala 39:30]
  wire  _T_296; // @[LZD.scala 39:27]
  wire  _T_297; // @[LZD.scala 39:25]
  wire [1:0] _T_298; // @[Cat.scala 29:58]
  wire [1:0] _T_299; // @[LZD.scala 44:32]
  wire  _T_300; // @[LZD.scala 39:14]
  wire  _T_301; // @[LZD.scala 39:21]
  wire  _T_302; // @[LZD.scala 39:30]
  wire  _T_303; // @[LZD.scala 39:27]
  wire  _T_304; // @[LZD.scala 39:25]
  wire [1:0] _T_305; // @[Cat.scala 29:58]
  wire  _T_306; // @[Shift.scala 12:21]
  wire  _T_307; // @[Shift.scala 12:21]
  wire  _T_308; // @[LZD.scala 49:16]
  wire  _T_309; // @[LZD.scala 49:27]
  wire  _T_310; // @[LZD.scala 49:25]
  wire  _T_311; // @[LZD.scala 49:47]
  wire  _T_312; // @[LZD.scala 49:59]
  wire  _T_313; // @[LZD.scala 49:35]
  wire [2:0] _T_315; // @[Cat.scala 29:58]
  wire [3:0] _T_316; // @[LZD.scala 44:32]
  wire [1:0] _T_317; // @[LZD.scala 43:32]
  wire  _T_318; // @[LZD.scala 39:14]
  wire  _T_319; // @[LZD.scala 39:21]
  wire  _T_320; // @[LZD.scala 39:30]
  wire  _T_321; // @[LZD.scala 39:27]
  wire  _T_322; // @[LZD.scala 39:25]
  wire [1:0] _T_323; // @[Cat.scala 29:58]
  wire [1:0] _T_324; // @[LZD.scala 44:32]
  wire  _T_325; // @[LZD.scala 39:14]
  wire  _T_326; // @[LZD.scala 39:21]
  wire  _T_327; // @[LZD.scala 39:30]
  wire  _T_328; // @[LZD.scala 39:27]
  wire  _T_329; // @[LZD.scala 39:25]
  wire [1:0] _T_330; // @[Cat.scala 29:58]
  wire  _T_331; // @[Shift.scala 12:21]
  wire  _T_332; // @[Shift.scala 12:21]
  wire  _T_333; // @[LZD.scala 49:16]
  wire  _T_334; // @[LZD.scala 49:27]
  wire  _T_335; // @[LZD.scala 49:25]
  wire  _T_336; // @[LZD.scala 49:47]
  wire  _T_337; // @[LZD.scala 49:59]
  wire  _T_338; // @[LZD.scala 49:35]
  wire [2:0] _T_340; // @[Cat.scala 29:58]
  wire  _T_341; // @[Shift.scala 12:21]
  wire  _T_342; // @[Shift.scala 12:21]
  wire  _T_343; // @[LZD.scala 49:16]
  wire  _T_344; // @[LZD.scala 49:27]
  wire  _T_345; // @[LZD.scala 49:25]
  wire [1:0] _T_346; // @[LZD.scala 49:47]
  wire [1:0] _T_347; // @[LZD.scala 49:59]
  wire [1:0] _T_348; // @[LZD.scala 49:35]
  wire [3:0] _T_350; // @[Cat.scala 29:58]
  wire [7:0] _T_351; // @[LZD.scala 44:32]
  wire [3:0] _T_352; // @[LZD.scala 43:32]
  wire [1:0] _T_353; // @[LZD.scala 43:32]
  wire  _T_354; // @[LZD.scala 39:14]
  wire  _T_355; // @[LZD.scala 39:21]
  wire  _T_356; // @[LZD.scala 39:30]
  wire  _T_357; // @[LZD.scala 39:27]
  wire  _T_358; // @[LZD.scala 39:25]
  wire [1:0] _T_359; // @[Cat.scala 29:58]
  wire [1:0] _T_360; // @[LZD.scala 44:32]
  wire  _T_361; // @[LZD.scala 39:14]
  wire  _T_362; // @[LZD.scala 39:21]
  wire  _T_363; // @[LZD.scala 39:30]
  wire  _T_364; // @[LZD.scala 39:27]
  wire  _T_365; // @[LZD.scala 39:25]
  wire [1:0] _T_366; // @[Cat.scala 29:58]
  wire  _T_367; // @[Shift.scala 12:21]
  wire  _T_368; // @[Shift.scala 12:21]
  wire  _T_369; // @[LZD.scala 49:16]
  wire  _T_370; // @[LZD.scala 49:27]
  wire  _T_371; // @[LZD.scala 49:25]
  wire  _T_372; // @[LZD.scala 49:47]
  wire  _T_373; // @[LZD.scala 49:59]
  wire  _T_374; // @[LZD.scala 49:35]
  wire [2:0] _T_376; // @[Cat.scala 29:58]
  wire [3:0] _T_377; // @[LZD.scala 44:32]
  wire [1:0] _T_378; // @[LZD.scala 43:32]
  wire  _T_379; // @[LZD.scala 39:14]
  wire  _T_380; // @[LZD.scala 39:21]
  wire  _T_381; // @[LZD.scala 39:30]
  wire  _T_382; // @[LZD.scala 39:27]
  wire  _T_383; // @[LZD.scala 39:25]
  wire [1:0] _T_384; // @[Cat.scala 29:58]
  wire [1:0] _T_385; // @[LZD.scala 44:32]
  wire  _T_386; // @[LZD.scala 39:14]
  wire  _T_387; // @[LZD.scala 39:21]
  wire  _T_388; // @[LZD.scala 39:30]
  wire  _T_389; // @[LZD.scala 39:27]
  wire  _T_390; // @[LZD.scala 39:25]
  wire [1:0] _T_391; // @[Cat.scala 29:58]
  wire  _T_392; // @[Shift.scala 12:21]
  wire  _T_393; // @[Shift.scala 12:21]
  wire  _T_394; // @[LZD.scala 49:16]
  wire  _T_395; // @[LZD.scala 49:27]
  wire  _T_396; // @[LZD.scala 49:25]
  wire  _T_397; // @[LZD.scala 49:47]
  wire  _T_398; // @[LZD.scala 49:59]
  wire  _T_399; // @[LZD.scala 49:35]
  wire [2:0] _T_401; // @[Cat.scala 29:58]
  wire  _T_402; // @[Shift.scala 12:21]
  wire  _T_403; // @[Shift.scala 12:21]
  wire  _T_404; // @[LZD.scala 49:16]
  wire  _T_405; // @[LZD.scala 49:27]
  wire  _T_406; // @[LZD.scala 49:25]
  wire [1:0] _T_407; // @[LZD.scala 49:47]
  wire [1:0] _T_408; // @[LZD.scala 49:59]
  wire [1:0] _T_409; // @[LZD.scala 49:35]
  wire [3:0] _T_411; // @[Cat.scala 29:58]
  wire  _T_412; // @[Shift.scala 12:21]
  wire  _T_413; // @[Shift.scala 12:21]
  wire  _T_414; // @[LZD.scala 49:16]
  wire  _T_415; // @[LZD.scala 49:27]
  wire  _T_416; // @[LZD.scala 49:25]
  wire [2:0] _T_417; // @[LZD.scala 49:47]
  wire [2:0] _T_418; // @[LZD.scala 49:59]
  wire [2:0] _T_419; // @[LZD.scala 49:35]
  wire [4:0] _T_421; // @[Cat.scala 29:58]
  wire [15:0] _T_422; // @[LZD.scala 44:32]
  wire [7:0] _T_423; // @[LZD.scala 43:32]
  wire [3:0] _T_424; // @[LZD.scala 43:32]
  wire [1:0] _T_425; // @[LZD.scala 43:32]
  wire  _T_426; // @[LZD.scala 39:14]
  wire  _T_427; // @[LZD.scala 39:21]
  wire  _T_428; // @[LZD.scala 39:30]
  wire  _T_429; // @[LZD.scala 39:27]
  wire  _T_430; // @[LZD.scala 39:25]
  wire [1:0] _T_431; // @[Cat.scala 29:58]
  wire [1:0] _T_432; // @[LZD.scala 44:32]
  wire  _T_433; // @[LZD.scala 39:14]
  wire  _T_434; // @[LZD.scala 39:21]
  wire  _T_435; // @[LZD.scala 39:30]
  wire  _T_436; // @[LZD.scala 39:27]
  wire  _T_437; // @[LZD.scala 39:25]
  wire [1:0] _T_438; // @[Cat.scala 29:58]
  wire  _T_439; // @[Shift.scala 12:21]
  wire  _T_440; // @[Shift.scala 12:21]
  wire  _T_441; // @[LZD.scala 49:16]
  wire  _T_442; // @[LZD.scala 49:27]
  wire  _T_443; // @[LZD.scala 49:25]
  wire  _T_444; // @[LZD.scala 49:47]
  wire  _T_445; // @[LZD.scala 49:59]
  wire  _T_446; // @[LZD.scala 49:35]
  wire [2:0] _T_448; // @[Cat.scala 29:58]
  wire [3:0] _T_449; // @[LZD.scala 44:32]
  wire [1:0] _T_450; // @[LZD.scala 43:32]
  wire  _T_451; // @[LZD.scala 39:14]
  wire  _T_452; // @[LZD.scala 39:21]
  wire  _T_453; // @[LZD.scala 39:30]
  wire  _T_454; // @[LZD.scala 39:27]
  wire  _T_455; // @[LZD.scala 39:25]
  wire [1:0] _T_456; // @[Cat.scala 29:58]
  wire [1:0] _T_457; // @[LZD.scala 44:32]
  wire  _T_458; // @[LZD.scala 39:14]
  wire  _T_459; // @[LZD.scala 39:21]
  wire  _T_460; // @[LZD.scala 39:30]
  wire  _T_461; // @[LZD.scala 39:27]
  wire  _T_462; // @[LZD.scala 39:25]
  wire [1:0] _T_463; // @[Cat.scala 29:58]
  wire  _T_464; // @[Shift.scala 12:21]
  wire  _T_465; // @[Shift.scala 12:21]
  wire  _T_466; // @[LZD.scala 49:16]
  wire  _T_467; // @[LZD.scala 49:27]
  wire  _T_468; // @[LZD.scala 49:25]
  wire  _T_469; // @[LZD.scala 49:47]
  wire  _T_470; // @[LZD.scala 49:59]
  wire  _T_471; // @[LZD.scala 49:35]
  wire [2:0] _T_473; // @[Cat.scala 29:58]
  wire  _T_474; // @[Shift.scala 12:21]
  wire  _T_475; // @[Shift.scala 12:21]
  wire  _T_476; // @[LZD.scala 49:16]
  wire  _T_477; // @[LZD.scala 49:27]
  wire  _T_478; // @[LZD.scala 49:25]
  wire [1:0] _T_479; // @[LZD.scala 49:47]
  wire [1:0] _T_480; // @[LZD.scala 49:59]
  wire [1:0] _T_481; // @[LZD.scala 49:35]
  wire [3:0] _T_483; // @[Cat.scala 29:58]
  wire [7:0] _T_484; // @[LZD.scala 44:32]
  wire [3:0] _T_485; // @[LZD.scala 43:32]
  wire [1:0] _T_486; // @[LZD.scala 43:32]
  wire  _T_487; // @[LZD.scala 39:14]
  wire  _T_488; // @[LZD.scala 39:21]
  wire  _T_489; // @[LZD.scala 39:30]
  wire  _T_490; // @[LZD.scala 39:27]
  wire  _T_491; // @[LZD.scala 39:25]
  wire [1:0] _T_492; // @[Cat.scala 29:58]
  wire [1:0] _T_493; // @[LZD.scala 44:32]
  wire  _T_494; // @[LZD.scala 39:14]
  wire  _T_495; // @[LZD.scala 39:21]
  wire  _T_496; // @[LZD.scala 39:30]
  wire  _T_497; // @[LZD.scala 39:27]
  wire  _T_498; // @[LZD.scala 39:25]
  wire [1:0] _T_499; // @[Cat.scala 29:58]
  wire  _T_500; // @[Shift.scala 12:21]
  wire  _T_501; // @[Shift.scala 12:21]
  wire  _T_502; // @[LZD.scala 49:16]
  wire  _T_503; // @[LZD.scala 49:27]
  wire  _T_504; // @[LZD.scala 49:25]
  wire  _T_505; // @[LZD.scala 49:47]
  wire  _T_506; // @[LZD.scala 49:59]
  wire  _T_507; // @[LZD.scala 49:35]
  wire [2:0] _T_509; // @[Cat.scala 29:58]
  wire [3:0] _T_510; // @[LZD.scala 44:32]
  wire [1:0] _T_511; // @[LZD.scala 43:32]
  wire  _T_512; // @[LZD.scala 39:14]
  wire  _T_513; // @[LZD.scala 39:21]
  wire  _T_514; // @[LZD.scala 39:30]
  wire  _T_515; // @[LZD.scala 39:27]
  wire  _T_516; // @[LZD.scala 39:25]
  wire [1:0] _T_517; // @[Cat.scala 29:58]
  wire [1:0] _T_518; // @[LZD.scala 44:32]
  wire  _T_519; // @[LZD.scala 39:14]
  wire  _T_520; // @[LZD.scala 39:21]
  wire  _T_521; // @[LZD.scala 39:30]
  wire  _T_522; // @[LZD.scala 39:27]
  wire  _T_523; // @[LZD.scala 39:25]
  wire [1:0] _T_524; // @[Cat.scala 29:58]
  wire  _T_525; // @[Shift.scala 12:21]
  wire  _T_526; // @[Shift.scala 12:21]
  wire  _T_527; // @[LZD.scala 49:16]
  wire  _T_528; // @[LZD.scala 49:27]
  wire  _T_529; // @[LZD.scala 49:25]
  wire  _T_530; // @[LZD.scala 49:47]
  wire  _T_531; // @[LZD.scala 49:59]
  wire  _T_532; // @[LZD.scala 49:35]
  wire [2:0] _T_534; // @[Cat.scala 29:58]
  wire  _T_535; // @[Shift.scala 12:21]
  wire  _T_536; // @[Shift.scala 12:21]
  wire  _T_537; // @[LZD.scala 49:16]
  wire  _T_538; // @[LZD.scala 49:27]
  wire  _T_539; // @[LZD.scala 49:25]
  wire [1:0] _T_540; // @[LZD.scala 49:47]
  wire [1:0] _T_541; // @[LZD.scala 49:59]
  wire [1:0] _T_542; // @[LZD.scala 49:35]
  wire [3:0] _T_544; // @[Cat.scala 29:58]
  wire  _T_545; // @[Shift.scala 12:21]
  wire  _T_546; // @[Shift.scala 12:21]
  wire  _T_547; // @[LZD.scala 49:16]
  wire  _T_548; // @[LZD.scala 49:27]
  wire  _T_549; // @[LZD.scala 49:25]
  wire [2:0] _T_550; // @[LZD.scala 49:47]
  wire [2:0] _T_551; // @[LZD.scala 49:59]
  wire [2:0] _T_552; // @[LZD.scala 49:35]
  wire [4:0] _T_554; // @[Cat.scala 29:58]
  wire  _T_555; // @[Shift.scala 12:21]
  wire  _T_556; // @[Shift.scala 12:21]
  wire  _T_557; // @[LZD.scala 49:16]
  wire  _T_558; // @[LZD.scala 49:27]
  wire  _T_559; // @[LZD.scala 49:25]
  wire [3:0] _T_560; // @[LZD.scala 49:47]
  wire [3:0] _T_561; // @[LZD.scala 49:59]
  wire [3:0] _T_562; // @[LZD.scala 49:35]
  wire [5:0] _T_564; // @[Cat.scala 29:58]
  wire  _T_565; // @[Shift.scala 12:21]
  wire  _T_566; // @[Shift.scala 12:21]
  wire  _T_567; // @[LZD.scala 49:16]
  wire  _T_568; // @[LZD.scala 49:27]
  wire  _T_569; // @[LZD.scala 49:25]
  wire [4:0] _T_570; // @[LZD.scala 49:47]
  wire [4:0] _T_571; // @[LZD.scala 49:59]
  wire [4:0] _T_572; // @[LZD.scala 49:35]
  wire [6:0] _T_574; // @[Cat.scala 29:58]
  wire [62:0] _T_575; // @[LZD.scala 44:32]
  wire [31:0] _T_576; // @[LZD.scala 43:32]
  wire [15:0] _T_577; // @[LZD.scala 43:32]
  wire [7:0] _T_578; // @[LZD.scala 43:32]
  wire [3:0] _T_579; // @[LZD.scala 43:32]
  wire [1:0] _T_580; // @[LZD.scala 43:32]
  wire  _T_581; // @[LZD.scala 39:14]
  wire  _T_582; // @[LZD.scala 39:21]
  wire  _T_583; // @[LZD.scala 39:30]
  wire  _T_584; // @[LZD.scala 39:27]
  wire  _T_585; // @[LZD.scala 39:25]
  wire [1:0] _T_586; // @[Cat.scala 29:58]
  wire [1:0] _T_587; // @[LZD.scala 44:32]
  wire  _T_588; // @[LZD.scala 39:14]
  wire  _T_589; // @[LZD.scala 39:21]
  wire  _T_590; // @[LZD.scala 39:30]
  wire  _T_591; // @[LZD.scala 39:27]
  wire  _T_592; // @[LZD.scala 39:25]
  wire [1:0] _T_593; // @[Cat.scala 29:58]
  wire  _T_594; // @[Shift.scala 12:21]
  wire  _T_595; // @[Shift.scala 12:21]
  wire  _T_596; // @[LZD.scala 49:16]
  wire  _T_597; // @[LZD.scala 49:27]
  wire  _T_598; // @[LZD.scala 49:25]
  wire  _T_599; // @[LZD.scala 49:47]
  wire  _T_600; // @[LZD.scala 49:59]
  wire  _T_601; // @[LZD.scala 49:35]
  wire [2:0] _T_603; // @[Cat.scala 29:58]
  wire [3:0] _T_604; // @[LZD.scala 44:32]
  wire [1:0] _T_605; // @[LZD.scala 43:32]
  wire  _T_606; // @[LZD.scala 39:14]
  wire  _T_607; // @[LZD.scala 39:21]
  wire  _T_608; // @[LZD.scala 39:30]
  wire  _T_609; // @[LZD.scala 39:27]
  wire  _T_610; // @[LZD.scala 39:25]
  wire [1:0] _T_611; // @[Cat.scala 29:58]
  wire [1:0] _T_612; // @[LZD.scala 44:32]
  wire  _T_613; // @[LZD.scala 39:14]
  wire  _T_614; // @[LZD.scala 39:21]
  wire  _T_615; // @[LZD.scala 39:30]
  wire  _T_616; // @[LZD.scala 39:27]
  wire  _T_617; // @[LZD.scala 39:25]
  wire [1:0] _T_618; // @[Cat.scala 29:58]
  wire  _T_619; // @[Shift.scala 12:21]
  wire  _T_620; // @[Shift.scala 12:21]
  wire  _T_621; // @[LZD.scala 49:16]
  wire  _T_622; // @[LZD.scala 49:27]
  wire  _T_623; // @[LZD.scala 49:25]
  wire  _T_624; // @[LZD.scala 49:47]
  wire  _T_625; // @[LZD.scala 49:59]
  wire  _T_626; // @[LZD.scala 49:35]
  wire [2:0] _T_628; // @[Cat.scala 29:58]
  wire  _T_629; // @[Shift.scala 12:21]
  wire  _T_630; // @[Shift.scala 12:21]
  wire  _T_631; // @[LZD.scala 49:16]
  wire  _T_632; // @[LZD.scala 49:27]
  wire  _T_633; // @[LZD.scala 49:25]
  wire [1:0] _T_634; // @[LZD.scala 49:47]
  wire [1:0] _T_635; // @[LZD.scala 49:59]
  wire [1:0] _T_636; // @[LZD.scala 49:35]
  wire [3:0] _T_638; // @[Cat.scala 29:58]
  wire [7:0] _T_639; // @[LZD.scala 44:32]
  wire [3:0] _T_640; // @[LZD.scala 43:32]
  wire [1:0] _T_641; // @[LZD.scala 43:32]
  wire  _T_642; // @[LZD.scala 39:14]
  wire  _T_643; // @[LZD.scala 39:21]
  wire  _T_644; // @[LZD.scala 39:30]
  wire  _T_645; // @[LZD.scala 39:27]
  wire  _T_646; // @[LZD.scala 39:25]
  wire [1:0] _T_647; // @[Cat.scala 29:58]
  wire [1:0] _T_648; // @[LZD.scala 44:32]
  wire  _T_649; // @[LZD.scala 39:14]
  wire  _T_650; // @[LZD.scala 39:21]
  wire  _T_651; // @[LZD.scala 39:30]
  wire  _T_652; // @[LZD.scala 39:27]
  wire  _T_653; // @[LZD.scala 39:25]
  wire [1:0] _T_654; // @[Cat.scala 29:58]
  wire  _T_655; // @[Shift.scala 12:21]
  wire  _T_656; // @[Shift.scala 12:21]
  wire  _T_657; // @[LZD.scala 49:16]
  wire  _T_658; // @[LZD.scala 49:27]
  wire  _T_659; // @[LZD.scala 49:25]
  wire  _T_660; // @[LZD.scala 49:47]
  wire  _T_661; // @[LZD.scala 49:59]
  wire  _T_662; // @[LZD.scala 49:35]
  wire [2:0] _T_664; // @[Cat.scala 29:58]
  wire [3:0] _T_665; // @[LZD.scala 44:32]
  wire [1:0] _T_666; // @[LZD.scala 43:32]
  wire  _T_667; // @[LZD.scala 39:14]
  wire  _T_668; // @[LZD.scala 39:21]
  wire  _T_669; // @[LZD.scala 39:30]
  wire  _T_670; // @[LZD.scala 39:27]
  wire  _T_671; // @[LZD.scala 39:25]
  wire [1:0] _T_672; // @[Cat.scala 29:58]
  wire [1:0] _T_673; // @[LZD.scala 44:32]
  wire  _T_674; // @[LZD.scala 39:14]
  wire  _T_675; // @[LZD.scala 39:21]
  wire  _T_676; // @[LZD.scala 39:30]
  wire  _T_677; // @[LZD.scala 39:27]
  wire  _T_678; // @[LZD.scala 39:25]
  wire [1:0] _T_679; // @[Cat.scala 29:58]
  wire  _T_680; // @[Shift.scala 12:21]
  wire  _T_681; // @[Shift.scala 12:21]
  wire  _T_682; // @[LZD.scala 49:16]
  wire  _T_683; // @[LZD.scala 49:27]
  wire  _T_684; // @[LZD.scala 49:25]
  wire  _T_685; // @[LZD.scala 49:47]
  wire  _T_686; // @[LZD.scala 49:59]
  wire  _T_687; // @[LZD.scala 49:35]
  wire [2:0] _T_689; // @[Cat.scala 29:58]
  wire  _T_690; // @[Shift.scala 12:21]
  wire  _T_691; // @[Shift.scala 12:21]
  wire  _T_692; // @[LZD.scala 49:16]
  wire  _T_693; // @[LZD.scala 49:27]
  wire  _T_694; // @[LZD.scala 49:25]
  wire [1:0] _T_695; // @[LZD.scala 49:47]
  wire [1:0] _T_696; // @[LZD.scala 49:59]
  wire [1:0] _T_697; // @[LZD.scala 49:35]
  wire [3:0] _T_699; // @[Cat.scala 29:58]
  wire  _T_700; // @[Shift.scala 12:21]
  wire  _T_701; // @[Shift.scala 12:21]
  wire  _T_702; // @[LZD.scala 49:16]
  wire  _T_703; // @[LZD.scala 49:27]
  wire  _T_704; // @[LZD.scala 49:25]
  wire [2:0] _T_705; // @[LZD.scala 49:47]
  wire [2:0] _T_706; // @[LZD.scala 49:59]
  wire [2:0] _T_707; // @[LZD.scala 49:35]
  wire [4:0] _T_709; // @[Cat.scala 29:58]
  wire [15:0] _T_710; // @[LZD.scala 44:32]
  wire [7:0] _T_711; // @[LZD.scala 43:32]
  wire [3:0] _T_712; // @[LZD.scala 43:32]
  wire [1:0] _T_713; // @[LZD.scala 43:32]
  wire  _T_714; // @[LZD.scala 39:14]
  wire  _T_715; // @[LZD.scala 39:21]
  wire  _T_716; // @[LZD.scala 39:30]
  wire  _T_717; // @[LZD.scala 39:27]
  wire  _T_718; // @[LZD.scala 39:25]
  wire [1:0] _T_719; // @[Cat.scala 29:58]
  wire [1:0] _T_720; // @[LZD.scala 44:32]
  wire  _T_721; // @[LZD.scala 39:14]
  wire  _T_722; // @[LZD.scala 39:21]
  wire  _T_723; // @[LZD.scala 39:30]
  wire  _T_724; // @[LZD.scala 39:27]
  wire  _T_725; // @[LZD.scala 39:25]
  wire [1:0] _T_726; // @[Cat.scala 29:58]
  wire  _T_727; // @[Shift.scala 12:21]
  wire  _T_728; // @[Shift.scala 12:21]
  wire  _T_729; // @[LZD.scala 49:16]
  wire  _T_730; // @[LZD.scala 49:27]
  wire  _T_731; // @[LZD.scala 49:25]
  wire  _T_732; // @[LZD.scala 49:47]
  wire  _T_733; // @[LZD.scala 49:59]
  wire  _T_734; // @[LZD.scala 49:35]
  wire [2:0] _T_736; // @[Cat.scala 29:58]
  wire [3:0] _T_737; // @[LZD.scala 44:32]
  wire [1:0] _T_738; // @[LZD.scala 43:32]
  wire  _T_739; // @[LZD.scala 39:14]
  wire  _T_740; // @[LZD.scala 39:21]
  wire  _T_741; // @[LZD.scala 39:30]
  wire  _T_742; // @[LZD.scala 39:27]
  wire  _T_743; // @[LZD.scala 39:25]
  wire [1:0] _T_744; // @[Cat.scala 29:58]
  wire [1:0] _T_745; // @[LZD.scala 44:32]
  wire  _T_746; // @[LZD.scala 39:14]
  wire  _T_747; // @[LZD.scala 39:21]
  wire  _T_748; // @[LZD.scala 39:30]
  wire  _T_749; // @[LZD.scala 39:27]
  wire  _T_750; // @[LZD.scala 39:25]
  wire [1:0] _T_751; // @[Cat.scala 29:58]
  wire  _T_752; // @[Shift.scala 12:21]
  wire  _T_753; // @[Shift.scala 12:21]
  wire  _T_754; // @[LZD.scala 49:16]
  wire  _T_755; // @[LZD.scala 49:27]
  wire  _T_756; // @[LZD.scala 49:25]
  wire  _T_757; // @[LZD.scala 49:47]
  wire  _T_758; // @[LZD.scala 49:59]
  wire  _T_759; // @[LZD.scala 49:35]
  wire [2:0] _T_761; // @[Cat.scala 29:58]
  wire  _T_762; // @[Shift.scala 12:21]
  wire  _T_763; // @[Shift.scala 12:21]
  wire  _T_764; // @[LZD.scala 49:16]
  wire  _T_765; // @[LZD.scala 49:27]
  wire  _T_766; // @[LZD.scala 49:25]
  wire [1:0] _T_767; // @[LZD.scala 49:47]
  wire [1:0] _T_768; // @[LZD.scala 49:59]
  wire [1:0] _T_769; // @[LZD.scala 49:35]
  wire [3:0] _T_771; // @[Cat.scala 29:58]
  wire [7:0] _T_772; // @[LZD.scala 44:32]
  wire [3:0] _T_773; // @[LZD.scala 43:32]
  wire [1:0] _T_774; // @[LZD.scala 43:32]
  wire  _T_775; // @[LZD.scala 39:14]
  wire  _T_776; // @[LZD.scala 39:21]
  wire  _T_777; // @[LZD.scala 39:30]
  wire  _T_778; // @[LZD.scala 39:27]
  wire  _T_779; // @[LZD.scala 39:25]
  wire [1:0] _T_780; // @[Cat.scala 29:58]
  wire [1:0] _T_781; // @[LZD.scala 44:32]
  wire  _T_782; // @[LZD.scala 39:14]
  wire  _T_783; // @[LZD.scala 39:21]
  wire  _T_784; // @[LZD.scala 39:30]
  wire  _T_785; // @[LZD.scala 39:27]
  wire  _T_786; // @[LZD.scala 39:25]
  wire [1:0] _T_787; // @[Cat.scala 29:58]
  wire  _T_788; // @[Shift.scala 12:21]
  wire  _T_789; // @[Shift.scala 12:21]
  wire  _T_790; // @[LZD.scala 49:16]
  wire  _T_791; // @[LZD.scala 49:27]
  wire  _T_792; // @[LZD.scala 49:25]
  wire  _T_793; // @[LZD.scala 49:47]
  wire  _T_794; // @[LZD.scala 49:59]
  wire  _T_795; // @[LZD.scala 49:35]
  wire [2:0] _T_797; // @[Cat.scala 29:58]
  wire [3:0] _T_798; // @[LZD.scala 44:32]
  wire [1:0] _T_799; // @[LZD.scala 43:32]
  wire  _T_800; // @[LZD.scala 39:14]
  wire  _T_801; // @[LZD.scala 39:21]
  wire  _T_802; // @[LZD.scala 39:30]
  wire  _T_803; // @[LZD.scala 39:27]
  wire  _T_804; // @[LZD.scala 39:25]
  wire [1:0] _T_805; // @[Cat.scala 29:58]
  wire [1:0] _T_806; // @[LZD.scala 44:32]
  wire  _T_807; // @[LZD.scala 39:14]
  wire  _T_808; // @[LZD.scala 39:21]
  wire  _T_809; // @[LZD.scala 39:30]
  wire  _T_810; // @[LZD.scala 39:27]
  wire  _T_811; // @[LZD.scala 39:25]
  wire [1:0] _T_812; // @[Cat.scala 29:58]
  wire  _T_813; // @[Shift.scala 12:21]
  wire  _T_814; // @[Shift.scala 12:21]
  wire  _T_815; // @[LZD.scala 49:16]
  wire  _T_816; // @[LZD.scala 49:27]
  wire  _T_817; // @[LZD.scala 49:25]
  wire  _T_818; // @[LZD.scala 49:47]
  wire  _T_819; // @[LZD.scala 49:59]
  wire  _T_820; // @[LZD.scala 49:35]
  wire [2:0] _T_822; // @[Cat.scala 29:58]
  wire  _T_823; // @[Shift.scala 12:21]
  wire  _T_824; // @[Shift.scala 12:21]
  wire  _T_825; // @[LZD.scala 49:16]
  wire  _T_826; // @[LZD.scala 49:27]
  wire  _T_827; // @[LZD.scala 49:25]
  wire [1:0] _T_828; // @[LZD.scala 49:47]
  wire [1:0] _T_829; // @[LZD.scala 49:59]
  wire [1:0] _T_830; // @[LZD.scala 49:35]
  wire [3:0] _T_832; // @[Cat.scala 29:58]
  wire  _T_833; // @[Shift.scala 12:21]
  wire  _T_834; // @[Shift.scala 12:21]
  wire  _T_835; // @[LZD.scala 49:16]
  wire  _T_836; // @[LZD.scala 49:27]
  wire  _T_837; // @[LZD.scala 49:25]
  wire [2:0] _T_838; // @[LZD.scala 49:47]
  wire [2:0] _T_839; // @[LZD.scala 49:59]
  wire [2:0] _T_840; // @[LZD.scala 49:35]
  wire [4:0] _T_842; // @[Cat.scala 29:58]
  wire  _T_843; // @[Shift.scala 12:21]
  wire  _T_844; // @[Shift.scala 12:21]
  wire  _T_845; // @[LZD.scala 49:16]
  wire  _T_846; // @[LZD.scala 49:27]
  wire  _T_847; // @[LZD.scala 49:25]
  wire [3:0] _T_848; // @[LZD.scala 49:47]
  wire [3:0] _T_849; // @[LZD.scala 49:59]
  wire [3:0] _T_850; // @[LZD.scala 49:35]
  wire [5:0] _T_852; // @[Cat.scala 29:58]
  wire [30:0] _T_853; // @[LZD.scala 44:32]
  wire [15:0] _T_854; // @[LZD.scala 43:32]
  wire [7:0] _T_855; // @[LZD.scala 43:32]
  wire [3:0] _T_856; // @[LZD.scala 43:32]
  wire [1:0] _T_857; // @[LZD.scala 43:32]
  wire  _T_858; // @[LZD.scala 39:14]
  wire  _T_859; // @[LZD.scala 39:21]
  wire  _T_860; // @[LZD.scala 39:30]
  wire  _T_861; // @[LZD.scala 39:27]
  wire  _T_862; // @[LZD.scala 39:25]
  wire [1:0] _T_863; // @[Cat.scala 29:58]
  wire [1:0] _T_864; // @[LZD.scala 44:32]
  wire  _T_865; // @[LZD.scala 39:14]
  wire  _T_866; // @[LZD.scala 39:21]
  wire  _T_867; // @[LZD.scala 39:30]
  wire  _T_868; // @[LZD.scala 39:27]
  wire  _T_869; // @[LZD.scala 39:25]
  wire [1:0] _T_870; // @[Cat.scala 29:58]
  wire  _T_871; // @[Shift.scala 12:21]
  wire  _T_872; // @[Shift.scala 12:21]
  wire  _T_873; // @[LZD.scala 49:16]
  wire  _T_874; // @[LZD.scala 49:27]
  wire  _T_875; // @[LZD.scala 49:25]
  wire  _T_876; // @[LZD.scala 49:47]
  wire  _T_877; // @[LZD.scala 49:59]
  wire  _T_878; // @[LZD.scala 49:35]
  wire [2:0] _T_880; // @[Cat.scala 29:58]
  wire [3:0] _T_881; // @[LZD.scala 44:32]
  wire [1:0] _T_882; // @[LZD.scala 43:32]
  wire  _T_883; // @[LZD.scala 39:14]
  wire  _T_884; // @[LZD.scala 39:21]
  wire  _T_885; // @[LZD.scala 39:30]
  wire  _T_886; // @[LZD.scala 39:27]
  wire  _T_887; // @[LZD.scala 39:25]
  wire [1:0] _T_888; // @[Cat.scala 29:58]
  wire [1:0] _T_889; // @[LZD.scala 44:32]
  wire  _T_890; // @[LZD.scala 39:14]
  wire  _T_891; // @[LZD.scala 39:21]
  wire  _T_892; // @[LZD.scala 39:30]
  wire  _T_893; // @[LZD.scala 39:27]
  wire  _T_894; // @[LZD.scala 39:25]
  wire [1:0] _T_895; // @[Cat.scala 29:58]
  wire  _T_896; // @[Shift.scala 12:21]
  wire  _T_897; // @[Shift.scala 12:21]
  wire  _T_898; // @[LZD.scala 49:16]
  wire  _T_899; // @[LZD.scala 49:27]
  wire  _T_900; // @[LZD.scala 49:25]
  wire  _T_901; // @[LZD.scala 49:47]
  wire  _T_902; // @[LZD.scala 49:59]
  wire  _T_903; // @[LZD.scala 49:35]
  wire [2:0] _T_905; // @[Cat.scala 29:58]
  wire  _T_906; // @[Shift.scala 12:21]
  wire  _T_907; // @[Shift.scala 12:21]
  wire  _T_908; // @[LZD.scala 49:16]
  wire  _T_909; // @[LZD.scala 49:27]
  wire  _T_910; // @[LZD.scala 49:25]
  wire [1:0] _T_911; // @[LZD.scala 49:47]
  wire [1:0] _T_912; // @[LZD.scala 49:59]
  wire [1:0] _T_913; // @[LZD.scala 49:35]
  wire [3:0] _T_915; // @[Cat.scala 29:58]
  wire [7:0] _T_916; // @[LZD.scala 44:32]
  wire [3:0] _T_917; // @[LZD.scala 43:32]
  wire [1:0] _T_918; // @[LZD.scala 43:32]
  wire  _T_919; // @[LZD.scala 39:14]
  wire  _T_920; // @[LZD.scala 39:21]
  wire  _T_921; // @[LZD.scala 39:30]
  wire  _T_922; // @[LZD.scala 39:27]
  wire  _T_923; // @[LZD.scala 39:25]
  wire [1:0] _T_924; // @[Cat.scala 29:58]
  wire [1:0] _T_925; // @[LZD.scala 44:32]
  wire  _T_926; // @[LZD.scala 39:14]
  wire  _T_927; // @[LZD.scala 39:21]
  wire  _T_928; // @[LZD.scala 39:30]
  wire  _T_929; // @[LZD.scala 39:27]
  wire  _T_930; // @[LZD.scala 39:25]
  wire [1:0] _T_931; // @[Cat.scala 29:58]
  wire  _T_932; // @[Shift.scala 12:21]
  wire  _T_933; // @[Shift.scala 12:21]
  wire  _T_934; // @[LZD.scala 49:16]
  wire  _T_935; // @[LZD.scala 49:27]
  wire  _T_936; // @[LZD.scala 49:25]
  wire  _T_937; // @[LZD.scala 49:47]
  wire  _T_938; // @[LZD.scala 49:59]
  wire  _T_939; // @[LZD.scala 49:35]
  wire [2:0] _T_941; // @[Cat.scala 29:58]
  wire [3:0] _T_942; // @[LZD.scala 44:32]
  wire [1:0] _T_943; // @[LZD.scala 43:32]
  wire  _T_944; // @[LZD.scala 39:14]
  wire  _T_945; // @[LZD.scala 39:21]
  wire  _T_946; // @[LZD.scala 39:30]
  wire  _T_947; // @[LZD.scala 39:27]
  wire  _T_948; // @[LZD.scala 39:25]
  wire [1:0] _T_949; // @[Cat.scala 29:58]
  wire [1:0] _T_950; // @[LZD.scala 44:32]
  wire  _T_951; // @[LZD.scala 39:14]
  wire  _T_952; // @[LZD.scala 39:21]
  wire  _T_953; // @[LZD.scala 39:30]
  wire  _T_954; // @[LZD.scala 39:27]
  wire  _T_955; // @[LZD.scala 39:25]
  wire [1:0] _T_956; // @[Cat.scala 29:58]
  wire  _T_957; // @[Shift.scala 12:21]
  wire  _T_958; // @[Shift.scala 12:21]
  wire  _T_959; // @[LZD.scala 49:16]
  wire  _T_960; // @[LZD.scala 49:27]
  wire  _T_961; // @[LZD.scala 49:25]
  wire  _T_962; // @[LZD.scala 49:47]
  wire  _T_963; // @[LZD.scala 49:59]
  wire  _T_964; // @[LZD.scala 49:35]
  wire [2:0] _T_966; // @[Cat.scala 29:58]
  wire  _T_967; // @[Shift.scala 12:21]
  wire  _T_968; // @[Shift.scala 12:21]
  wire  _T_969; // @[LZD.scala 49:16]
  wire  _T_970; // @[LZD.scala 49:27]
  wire  _T_971; // @[LZD.scala 49:25]
  wire [1:0] _T_972; // @[LZD.scala 49:47]
  wire [1:0] _T_973; // @[LZD.scala 49:59]
  wire [1:0] _T_974; // @[LZD.scala 49:35]
  wire [3:0] _T_976; // @[Cat.scala 29:58]
  wire  _T_977; // @[Shift.scala 12:21]
  wire  _T_978; // @[Shift.scala 12:21]
  wire  _T_979; // @[LZD.scala 49:16]
  wire  _T_980; // @[LZD.scala 49:27]
  wire  _T_981; // @[LZD.scala 49:25]
  wire [2:0] _T_982; // @[LZD.scala 49:47]
  wire [2:0] _T_983; // @[LZD.scala 49:59]
  wire [2:0] _T_984; // @[LZD.scala 49:35]
  wire [4:0] _T_986; // @[Cat.scala 29:58]
  wire [14:0] _T_987; // @[LZD.scala 44:32]
  wire [7:0] _T_988; // @[LZD.scala 43:32]
  wire [3:0] _T_989; // @[LZD.scala 43:32]
  wire [1:0] _T_990; // @[LZD.scala 43:32]
  wire  _T_991; // @[LZD.scala 39:14]
  wire  _T_992; // @[LZD.scala 39:21]
  wire  _T_993; // @[LZD.scala 39:30]
  wire  _T_994; // @[LZD.scala 39:27]
  wire  _T_995; // @[LZD.scala 39:25]
  wire [1:0] _T_996; // @[Cat.scala 29:58]
  wire [1:0] _T_997; // @[LZD.scala 44:32]
  wire  _T_998; // @[LZD.scala 39:14]
  wire  _T_999; // @[LZD.scala 39:21]
  wire  _T_1000; // @[LZD.scala 39:30]
  wire  _T_1001; // @[LZD.scala 39:27]
  wire  _T_1002; // @[LZD.scala 39:25]
  wire [1:0] _T_1003; // @[Cat.scala 29:58]
  wire  _T_1004; // @[Shift.scala 12:21]
  wire  _T_1005; // @[Shift.scala 12:21]
  wire  _T_1006; // @[LZD.scala 49:16]
  wire  _T_1007; // @[LZD.scala 49:27]
  wire  _T_1008; // @[LZD.scala 49:25]
  wire  _T_1009; // @[LZD.scala 49:47]
  wire  _T_1010; // @[LZD.scala 49:59]
  wire  _T_1011; // @[LZD.scala 49:35]
  wire [2:0] _T_1013; // @[Cat.scala 29:58]
  wire [3:0] _T_1014; // @[LZD.scala 44:32]
  wire [1:0] _T_1015; // @[LZD.scala 43:32]
  wire  _T_1016; // @[LZD.scala 39:14]
  wire  _T_1017; // @[LZD.scala 39:21]
  wire  _T_1018; // @[LZD.scala 39:30]
  wire  _T_1019; // @[LZD.scala 39:27]
  wire  _T_1020; // @[LZD.scala 39:25]
  wire [1:0] _T_1021; // @[Cat.scala 29:58]
  wire [1:0] _T_1022; // @[LZD.scala 44:32]
  wire  _T_1023; // @[LZD.scala 39:14]
  wire  _T_1024; // @[LZD.scala 39:21]
  wire  _T_1025; // @[LZD.scala 39:30]
  wire  _T_1026; // @[LZD.scala 39:27]
  wire  _T_1027; // @[LZD.scala 39:25]
  wire [1:0] _T_1028; // @[Cat.scala 29:58]
  wire  _T_1029; // @[Shift.scala 12:21]
  wire  _T_1030; // @[Shift.scala 12:21]
  wire  _T_1031; // @[LZD.scala 49:16]
  wire  _T_1032; // @[LZD.scala 49:27]
  wire  _T_1033; // @[LZD.scala 49:25]
  wire  _T_1034; // @[LZD.scala 49:47]
  wire  _T_1035; // @[LZD.scala 49:59]
  wire  _T_1036; // @[LZD.scala 49:35]
  wire [2:0] _T_1038; // @[Cat.scala 29:58]
  wire  _T_1039; // @[Shift.scala 12:21]
  wire  _T_1040; // @[Shift.scala 12:21]
  wire  _T_1041; // @[LZD.scala 49:16]
  wire  _T_1042; // @[LZD.scala 49:27]
  wire  _T_1043; // @[LZD.scala 49:25]
  wire [1:0] _T_1044; // @[LZD.scala 49:47]
  wire [1:0] _T_1045; // @[LZD.scala 49:59]
  wire [1:0] _T_1046; // @[LZD.scala 49:35]
  wire [3:0] _T_1048; // @[Cat.scala 29:58]
  wire [6:0] _T_1049; // @[LZD.scala 44:32]
  wire [3:0] _T_1050; // @[LZD.scala 43:32]
  wire [1:0] _T_1051; // @[LZD.scala 43:32]
  wire  _T_1052; // @[LZD.scala 39:14]
  wire  _T_1053; // @[LZD.scala 39:21]
  wire  _T_1054; // @[LZD.scala 39:30]
  wire  _T_1055; // @[LZD.scala 39:27]
  wire  _T_1056; // @[LZD.scala 39:25]
  wire [1:0] _T_1057; // @[Cat.scala 29:58]
  wire [1:0] _T_1058; // @[LZD.scala 44:32]
  wire  _T_1059; // @[LZD.scala 39:14]
  wire  _T_1060; // @[LZD.scala 39:21]
  wire  _T_1061; // @[LZD.scala 39:30]
  wire  _T_1062; // @[LZD.scala 39:27]
  wire  _T_1063; // @[LZD.scala 39:25]
  wire [1:0] _T_1064; // @[Cat.scala 29:58]
  wire  _T_1065; // @[Shift.scala 12:21]
  wire  _T_1066; // @[Shift.scala 12:21]
  wire  _T_1067; // @[LZD.scala 49:16]
  wire  _T_1068; // @[LZD.scala 49:27]
  wire  _T_1069; // @[LZD.scala 49:25]
  wire  _T_1070; // @[LZD.scala 49:47]
  wire  _T_1071; // @[LZD.scala 49:59]
  wire  _T_1072; // @[LZD.scala 49:35]
  wire [2:0] _T_1074; // @[Cat.scala 29:58]
  wire [2:0] _T_1075; // @[LZD.scala 44:32]
  wire [1:0] _T_1076; // @[LZD.scala 43:32]
  wire  _T_1077; // @[LZD.scala 39:14]
  wire  _T_1078; // @[LZD.scala 39:21]
  wire  _T_1079; // @[LZD.scala 39:30]
  wire  _T_1080; // @[LZD.scala 39:27]
  wire  _T_1081; // @[LZD.scala 39:25]
  wire [1:0] _T_1082; // @[Cat.scala 29:58]
  wire  _T_1083; // @[LZD.scala 44:32]
  wire  _T_1085; // @[Shift.scala 12:21]
  wire  _T_1087; // @[LZD.scala 55:32]
  wire  _T_1088; // @[LZD.scala 55:20]
  wire [1:0] _T_1089; // @[Cat.scala 29:58]
  wire  _T_1090; // @[Shift.scala 12:21]
  wire [1:0] _T_1092; // @[LZD.scala 55:32]
  wire [1:0] _T_1093; // @[LZD.scala 55:20]
  wire [2:0] _T_1094; // @[Cat.scala 29:58]
  wire  _T_1095; // @[Shift.scala 12:21]
  wire [2:0] _T_1097; // @[LZD.scala 55:32]
  wire [2:0] _T_1098; // @[LZD.scala 55:20]
  wire [3:0] _T_1099; // @[Cat.scala 29:58]
  wire  _T_1100; // @[Shift.scala 12:21]
  wire [3:0] _T_1102; // @[LZD.scala 55:32]
  wire [3:0] _T_1103; // @[LZD.scala 55:20]
  wire [4:0] _T_1104; // @[Cat.scala 29:58]
  wire  _T_1105; // @[Shift.scala 12:21]
  wire [4:0] _T_1107; // @[LZD.scala 55:32]
  wire [4:0] _T_1108; // @[LZD.scala 55:20]
  wire [5:0] _T_1109; // @[Cat.scala 29:58]
  wire  _T_1110; // @[Shift.scala 12:21]
  wire [5:0] _T_1112; // @[LZD.scala 55:32]
  wire [5:0] _T_1113; // @[LZD.scala 55:20]
  wire [7:0] scaleBias; // @[Cat.scala 29:58]
  wire [7:0] _T_1114; // @[QuireToPosit.scala 61:53]
  wire [8:0] _GEN_2; // @[QuireToPosit.scala 61:41]
  wire [8:0] _T_1116; // @[QuireToPosit.scala 61:41]
  wire [8:0] realScale; // @[QuireToPosit.scala 61:41]
  wire  underflow; // @[QuireToPosit.scala 62:41]
  wire  overflow; // @[QuireToPosit.scala 63:35]
  wire [8:0] _T_1117; // @[Mux.scala 87:16]
  wire [8:0] _T_1118; // @[Mux.scala 87:16]
  wire  _T_1119; // @[Abs.scala 10:21]
  wire [8:0] _T_1121; // @[Bitwise.scala 71:12]
  wire [8:0] _T_1122; // @[Abs.scala 10:31]
  wire [8:0] _T_1123; // @[Abs.scala 10:26]
  wire [8:0] _GEN_3; // @[Abs.scala 10:39]
  wire [8:0] absRealScale; // @[Abs.scala 10:39]
  wire  _T_1126; // @[Shift.scala 16:24]
  wire [6:0] _T_1127; // @[Shift.scala 17:37]
  wire  _T_1128; // @[Shift.scala 12:21]
  wire [63:0] _T_1129; // @[Shift.scala 64:52]
  wire [127:0] _T_1131; // @[Cat.scala 29:58]
  wire [127:0] _T_1132; // @[Shift.scala 64:27]
  wire [5:0] _T_1133; // @[Shift.scala 66:70]
  wire  _T_1134; // @[Shift.scala 12:21]
  wire [95:0] _T_1135; // @[Shift.scala 64:52]
  wire [127:0] _T_1137; // @[Cat.scala 29:58]
  wire [127:0] _T_1138; // @[Shift.scala 64:27]
  wire [4:0] _T_1139; // @[Shift.scala 66:70]
  wire  _T_1140; // @[Shift.scala 12:21]
  wire [111:0] _T_1141; // @[Shift.scala 64:52]
  wire [127:0] _T_1143; // @[Cat.scala 29:58]
  wire [127:0] _T_1144; // @[Shift.scala 64:27]
  wire [3:0] _T_1145; // @[Shift.scala 66:70]
  wire  _T_1146; // @[Shift.scala 12:21]
  wire [119:0] _T_1147; // @[Shift.scala 64:52]
  wire [127:0] _T_1149; // @[Cat.scala 29:58]
  wire [127:0] _T_1150; // @[Shift.scala 64:27]
  wire [2:0] _T_1151; // @[Shift.scala 66:70]
  wire  _T_1152; // @[Shift.scala 12:21]
  wire [123:0] _T_1153; // @[Shift.scala 64:52]
  wire [127:0] _T_1155; // @[Cat.scala 29:58]
  wire [127:0] _T_1156; // @[Shift.scala 64:27]
  wire [1:0] _T_1157; // @[Shift.scala 66:70]
  wire  _T_1158; // @[Shift.scala 12:21]
  wire [125:0] _T_1159; // @[Shift.scala 64:52]
  wire [127:0] _T_1161; // @[Cat.scala 29:58]
  wire [127:0] _T_1162; // @[Shift.scala 64:27]
  wire  _T_1163; // @[Shift.scala 66:70]
  wire [126:0] _T_1165; // @[Shift.scala 64:52]
  wire [127:0] _T_1166; // @[Cat.scala 29:58]
  wire [127:0] _T_1167; // @[Shift.scala 64:27]
  wire [127:0] quireLeftShift; // @[Shift.scala 16:10]
  wire [63:0] _T_1172; // @[Shift.scala 77:66]
  wire [127:0] _T_1173; // @[Cat.scala 29:58]
  wire [127:0] _T_1174; // @[Shift.scala 77:22]
  wire [95:0] _T_1178; // @[Shift.scala 77:66]
  wire [127:0] _T_1179; // @[Cat.scala 29:58]
  wire [127:0] _T_1180; // @[Shift.scala 77:22]
  wire [111:0] _T_1184; // @[Shift.scala 77:66]
  wire [127:0] _T_1185; // @[Cat.scala 29:58]
  wire [127:0] _T_1186; // @[Shift.scala 77:22]
  wire [119:0] _T_1190; // @[Shift.scala 77:66]
  wire [127:0] _T_1191; // @[Cat.scala 29:58]
  wire [127:0] _T_1192; // @[Shift.scala 77:22]
  wire [123:0] _T_1196; // @[Shift.scala 77:66]
  wire [127:0] _T_1197; // @[Cat.scala 29:58]
  wire [127:0] _T_1198; // @[Shift.scala 77:22]
  wire [125:0] _T_1202; // @[Shift.scala 77:66]
  wire [127:0] _T_1203; // @[Cat.scala 29:58]
  wire [127:0] _T_1204; // @[Shift.scala 77:22]
  wire [126:0] _T_1207; // @[Shift.scala 77:66]
  wire [127:0] _T_1208; // @[Cat.scala 29:58]
  wire [127:0] _T_1209; // @[Shift.scala 77:22]
  wire [127:0] quireRightShift; // @[Shift.scala 27:10]
  wire [4:0] _T_1211; // @[QuireToPosit.scala 89:49]
  wire [42:0] _T_1212; // @[QuireToPosit.scala 90:127]
  wire  _T_1213; // @[QuireToPosit.scala 90:154]
  wire [5:0] realFGRSTmp1; // @[Cat.scala 29:58]
  wire [4:0] _T_1214; // @[QuireToPosit.scala 91:50]
  wire [42:0] _T_1215; // @[QuireToPosit.scala 92:128]
  wire  _T_1216; // @[QuireToPosit.scala 92:155]
  wire [5:0] realFGRSTmp2; // @[Cat.scala 29:58]
  wire [5:0] realFGRS; // @[QuireToPosit.scala 93:34]
  wire [2:0] outRawFloat_fraction; // @[QuireToPosit.scala 95:46]
  wire [2:0] outRawFloat_grs; // @[QuireToPosit.scala 96:46]
  wire [5:0] _GEN_4; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire [5:0] outRawFloat_scale; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  wire [1:0] _T_1221; // @[convert.scala 46:61]
  wire [1:0] _T_1222; // @[convert.scala 46:52]
  wire [1:0] _T_1224; // @[convert.scala 46:42]
  wire [3:0] _T_1225; // @[convert.scala 48:34]
  wire  _T_1226; // @[convert.scala 49:36]
  wire [3:0] _T_1228; // @[convert.scala 50:36]
  wire [3:0] _T_1229; // @[convert.scala 50:36]
  wire [3:0] _T_1230; // @[convert.scala 50:28]
  wire  _T_1231; // @[convert.scala 51:31]
  wire  _T_1232; // @[convert.scala 52:43]
  wire [9:0] _T_1236; // @[Cat.scala 29:58]
  wire [3:0] _T_1237; // @[Shift.scala 39:17]
  wire  _T_1238; // @[Shift.scala 39:24]
  wire [1:0] _T_1240; // @[Shift.scala 90:30]
  wire [7:0] _T_1241; // @[Shift.scala 90:48]
  wire  _T_1242; // @[Shift.scala 90:57]
  wire [1:0] _GEN_5; // @[Shift.scala 90:39]
  wire [1:0] _T_1243; // @[Shift.scala 90:39]
  wire  _T_1244; // @[Shift.scala 12:21]
  wire  _T_1245; // @[Shift.scala 12:21]
  wire [7:0] _T_1247; // @[Bitwise.scala 71:12]
  wire [9:0] _T_1248; // @[Cat.scala 29:58]
  wire [9:0] _T_1249; // @[Shift.scala 91:22]
  wire [2:0] _T_1250; // @[Shift.scala 92:77]
  wire [5:0] _T_1251; // @[Shift.scala 90:30]
  wire [3:0] _T_1252; // @[Shift.scala 90:48]
  wire  _T_1253; // @[Shift.scala 90:57]
  wire [5:0] _GEN_6; // @[Shift.scala 90:39]
  wire [5:0] _T_1254; // @[Shift.scala 90:39]
  wire  _T_1255; // @[Shift.scala 12:21]
  wire  _T_1256; // @[Shift.scala 12:21]
  wire [3:0] _T_1258; // @[Bitwise.scala 71:12]
  wire [9:0] _T_1259; // @[Cat.scala 29:58]
  wire [9:0] _T_1260; // @[Shift.scala 91:22]
  wire [1:0] _T_1261; // @[Shift.scala 92:77]
  wire [7:0] _T_1262; // @[Shift.scala 90:30]
  wire [1:0] _T_1263; // @[Shift.scala 90:48]
  wire  _T_1264; // @[Shift.scala 90:57]
  wire [7:0] _GEN_7; // @[Shift.scala 90:39]
  wire [7:0] _T_1265; // @[Shift.scala 90:39]
  wire  _T_1266; // @[Shift.scala 12:21]
  wire  _T_1267; // @[Shift.scala 12:21]
  wire [1:0] _T_1269; // @[Bitwise.scala 71:12]
  wire [9:0] _T_1270; // @[Cat.scala 29:58]
  wire [9:0] _T_1271; // @[Shift.scala 91:22]
  wire  _T_1272; // @[Shift.scala 92:77]
  wire [8:0] _T_1273; // @[Shift.scala 90:30]
  wire  _T_1274; // @[Shift.scala 90:48]
  wire [8:0] _GEN_8; // @[Shift.scala 90:39]
  wire [8:0] _T_1276; // @[Shift.scala 90:39]
  wire  _T_1278; // @[Shift.scala 12:21]
  wire [9:0] _T_1279; // @[Cat.scala 29:58]
  wire [9:0] _T_1280; // @[Shift.scala 91:22]
  wire [9:0] _T_1283; // @[Bitwise.scala 71:12]
  wire [9:0] _T_1284; // @[Shift.scala 39:10]
  wire  _T_1285; // @[convert.scala 55:31]
  wire  _T_1286; // @[convert.scala 56:31]
  wire  _T_1287; // @[convert.scala 57:31]
  wire  _T_1288; // @[convert.scala 58:31]
  wire [6:0] _T_1289; // @[convert.scala 59:69]
  wire  _T_1290; // @[convert.scala 59:81]
  wire  _T_1291; // @[convert.scala 59:50]
  wire  _T_1293; // @[convert.scala 60:81]
  wire  _T_1294; // @[convert.scala 61:44]
  wire  _T_1295; // @[convert.scala 61:52]
  wire  _T_1296; // @[convert.scala 61:36]
  wire  _T_1297; // @[convert.scala 62:63]
  wire  _T_1298; // @[convert.scala 62:103]
  wire  _T_1299; // @[convert.scala 62:60]
  wire [6:0] _GEN_9; // @[convert.scala 63:56]
  wire [6:0] _T_1302; // @[convert.scala 63:56]
  wire [7:0] _T_1303; // @[Cat.scala 29:58]
  reg  _T_1307; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1311; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  assign _T = io_quireIn[126:0]; // @[QuireToPosit.scala 47:43]
  assign _T_1 = _T != 127'h0; // @[QuireToPosit.scala 47:47]
  assign tailIsZero = ~ _T_1; // @[QuireToPosit.scala 47:27]
  assign _T_2 = io_quireIn[127:127]; // @[QuireToPosit.scala 49:45]
  assign outRawFloat_isNaR = _T_2 & tailIsZero; // @[QuireToPosit.scala 49:49]
  assign _T_5 = ~ _T_2; // @[QuireToPosit.scala 50:31]
  assign outRawFloat_isZero = _T_5 & tailIsZero; // @[QuireToPosit.scala 50:51]
  assign _T_8 = io_quireIn[127:1]; // @[QuireToPosit.scala 58:41]
  assign _T_9 = io_quireIn[126:0]; // @[QuireToPosit.scala 58:68]
  assign quireXOR = _T_8 ^ _T_9; // @[QuireToPosit.scala 58:56]
  assign _T_10 = quireXOR[126:63]; // @[LZD.scala 43:32]
  assign _T_11 = _T_10[63:32]; // @[LZD.scala 43:32]
  assign _T_12 = _T_11[31:16]; // @[LZD.scala 43:32]
  assign _T_13 = _T_12[15:8]; // @[LZD.scala 43:32]
  assign _T_14 = _T_13[7:4]; // @[LZD.scala 43:32]
  assign _T_15 = _T_14[3:2]; // @[LZD.scala 43:32]
  assign _T_16 = _T_15 != 2'h0; // @[LZD.scala 39:14]
  assign _T_17 = _T_15[1]; // @[LZD.scala 39:21]
  assign _T_18 = _T_15[0]; // @[LZD.scala 39:30]
  assign _T_19 = ~ _T_18; // @[LZD.scala 39:27]
  assign _T_20 = _T_17 | _T_19; // @[LZD.scala 39:25]
  assign _T_21 = {_T_16,_T_20}; // @[Cat.scala 29:58]
  assign _T_22 = _T_14[1:0]; // @[LZD.scala 44:32]
  assign _T_23 = _T_22 != 2'h0; // @[LZD.scala 39:14]
  assign _T_24 = _T_22[1]; // @[LZD.scala 39:21]
  assign _T_25 = _T_22[0]; // @[LZD.scala 39:30]
  assign _T_26 = ~ _T_25; // @[LZD.scala 39:27]
  assign _T_27 = _T_24 | _T_26; // @[LZD.scala 39:25]
  assign _T_28 = {_T_23,_T_27}; // @[Cat.scala 29:58]
  assign _T_29 = _T_21[1]; // @[Shift.scala 12:21]
  assign _T_30 = _T_28[1]; // @[Shift.scala 12:21]
  assign _T_31 = _T_29 | _T_30; // @[LZD.scala 49:16]
  assign _T_32 = ~ _T_30; // @[LZD.scala 49:27]
  assign _T_33 = _T_29 | _T_32; // @[LZD.scala 49:25]
  assign _T_34 = _T_21[0:0]; // @[LZD.scala 49:47]
  assign _T_35 = _T_28[0:0]; // @[LZD.scala 49:59]
  assign _T_36 = _T_29 ? _T_34 : _T_35; // @[LZD.scala 49:35]
  assign _T_38 = {_T_31,_T_33,_T_36}; // @[Cat.scala 29:58]
  assign _T_39 = _T_13[3:0]; // @[LZD.scala 44:32]
  assign _T_40 = _T_39[3:2]; // @[LZD.scala 43:32]
  assign _T_41 = _T_40 != 2'h0; // @[LZD.scala 39:14]
  assign _T_42 = _T_40[1]; // @[LZD.scala 39:21]
  assign _T_43 = _T_40[0]; // @[LZD.scala 39:30]
  assign _T_44 = ~ _T_43; // @[LZD.scala 39:27]
  assign _T_45 = _T_42 | _T_44; // @[LZD.scala 39:25]
  assign _T_46 = {_T_41,_T_45}; // @[Cat.scala 29:58]
  assign _T_47 = _T_39[1:0]; // @[LZD.scala 44:32]
  assign _T_48 = _T_47 != 2'h0; // @[LZD.scala 39:14]
  assign _T_49 = _T_47[1]; // @[LZD.scala 39:21]
  assign _T_50 = _T_47[0]; // @[LZD.scala 39:30]
  assign _T_51 = ~ _T_50; // @[LZD.scala 39:27]
  assign _T_52 = _T_49 | _T_51; // @[LZD.scala 39:25]
  assign _T_53 = {_T_48,_T_52}; // @[Cat.scala 29:58]
  assign _T_54 = _T_46[1]; // @[Shift.scala 12:21]
  assign _T_55 = _T_53[1]; // @[Shift.scala 12:21]
  assign _T_56 = _T_54 | _T_55; // @[LZD.scala 49:16]
  assign _T_57 = ~ _T_55; // @[LZD.scala 49:27]
  assign _T_58 = _T_54 | _T_57; // @[LZD.scala 49:25]
  assign _T_59 = _T_46[0:0]; // @[LZD.scala 49:47]
  assign _T_60 = _T_53[0:0]; // @[LZD.scala 49:59]
  assign _T_61 = _T_54 ? _T_59 : _T_60; // @[LZD.scala 49:35]
  assign _T_63 = {_T_56,_T_58,_T_61}; // @[Cat.scala 29:58]
  assign _T_64 = _T_38[2]; // @[Shift.scala 12:21]
  assign _T_65 = _T_63[2]; // @[Shift.scala 12:21]
  assign _T_66 = _T_64 | _T_65; // @[LZD.scala 49:16]
  assign _T_67 = ~ _T_65; // @[LZD.scala 49:27]
  assign _T_68 = _T_64 | _T_67; // @[LZD.scala 49:25]
  assign _T_69 = _T_38[1:0]; // @[LZD.scala 49:47]
  assign _T_70 = _T_63[1:0]; // @[LZD.scala 49:59]
  assign _T_71 = _T_64 ? _T_69 : _T_70; // @[LZD.scala 49:35]
  assign _T_73 = {_T_66,_T_68,_T_71}; // @[Cat.scala 29:58]
  assign _T_74 = _T_12[7:0]; // @[LZD.scala 44:32]
  assign _T_75 = _T_74[7:4]; // @[LZD.scala 43:32]
  assign _T_76 = _T_75[3:2]; // @[LZD.scala 43:32]
  assign _T_77 = _T_76 != 2'h0; // @[LZD.scala 39:14]
  assign _T_78 = _T_76[1]; // @[LZD.scala 39:21]
  assign _T_79 = _T_76[0]; // @[LZD.scala 39:30]
  assign _T_80 = ~ _T_79; // @[LZD.scala 39:27]
  assign _T_81 = _T_78 | _T_80; // @[LZD.scala 39:25]
  assign _T_82 = {_T_77,_T_81}; // @[Cat.scala 29:58]
  assign _T_83 = _T_75[1:0]; // @[LZD.scala 44:32]
  assign _T_84 = _T_83 != 2'h0; // @[LZD.scala 39:14]
  assign _T_85 = _T_83[1]; // @[LZD.scala 39:21]
  assign _T_86 = _T_83[0]; // @[LZD.scala 39:30]
  assign _T_87 = ~ _T_86; // @[LZD.scala 39:27]
  assign _T_88 = _T_85 | _T_87; // @[LZD.scala 39:25]
  assign _T_89 = {_T_84,_T_88}; // @[Cat.scala 29:58]
  assign _T_90 = _T_82[1]; // @[Shift.scala 12:21]
  assign _T_91 = _T_89[1]; // @[Shift.scala 12:21]
  assign _T_92 = _T_90 | _T_91; // @[LZD.scala 49:16]
  assign _T_93 = ~ _T_91; // @[LZD.scala 49:27]
  assign _T_94 = _T_90 | _T_93; // @[LZD.scala 49:25]
  assign _T_95 = _T_82[0:0]; // @[LZD.scala 49:47]
  assign _T_96 = _T_89[0:0]; // @[LZD.scala 49:59]
  assign _T_97 = _T_90 ? _T_95 : _T_96; // @[LZD.scala 49:35]
  assign _T_99 = {_T_92,_T_94,_T_97}; // @[Cat.scala 29:58]
  assign _T_100 = _T_74[3:0]; // @[LZD.scala 44:32]
  assign _T_101 = _T_100[3:2]; // @[LZD.scala 43:32]
  assign _T_102 = _T_101 != 2'h0; // @[LZD.scala 39:14]
  assign _T_103 = _T_101[1]; // @[LZD.scala 39:21]
  assign _T_104 = _T_101[0]; // @[LZD.scala 39:30]
  assign _T_105 = ~ _T_104; // @[LZD.scala 39:27]
  assign _T_106 = _T_103 | _T_105; // @[LZD.scala 39:25]
  assign _T_107 = {_T_102,_T_106}; // @[Cat.scala 29:58]
  assign _T_108 = _T_100[1:0]; // @[LZD.scala 44:32]
  assign _T_109 = _T_108 != 2'h0; // @[LZD.scala 39:14]
  assign _T_110 = _T_108[1]; // @[LZD.scala 39:21]
  assign _T_111 = _T_108[0]; // @[LZD.scala 39:30]
  assign _T_112 = ~ _T_111; // @[LZD.scala 39:27]
  assign _T_113 = _T_110 | _T_112; // @[LZD.scala 39:25]
  assign _T_114 = {_T_109,_T_113}; // @[Cat.scala 29:58]
  assign _T_115 = _T_107[1]; // @[Shift.scala 12:21]
  assign _T_116 = _T_114[1]; // @[Shift.scala 12:21]
  assign _T_117 = _T_115 | _T_116; // @[LZD.scala 49:16]
  assign _T_118 = ~ _T_116; // @[LZD.scala 49:27]
  assign _T_119 = _T_115 | _T_118; // @[LZD.scala 49:25]
  assign _T_120 = _T_107[0:0]; // @[LZD.scala 49:47]
  assign _T_121 = _T_114[0:0]; // @[LZD.scala 49:59]
  assign _T_122 = _T_115 ? _T_120 : _T_121; // @[LZD.scala 49:35]
  assign _T_124 = {_T_117,_T_119,_T_122}; // @[Cat.scala 29:58]
  assign _T_125 = _T_99[2]; // @[Shift.scala 12:21]
  assign _T_126 = _T_124[2]; // @[Shift.scala 12:21]
  assign _T_127 = _T_125 | _T_126; // @[LZD.scala 49:16]
  assign _T_128 = ~ _T_126; // @[LZD.scala 49:27]
  assign _T_129 = _T_125 | _T_128; // @[LZD.scala 49:25]
  assign _T_130 = _T_99[1:0]; // @[LZD.scala 49:47]
  assign _T_131 = _T_124[1:0]; // @[LZD.scala 49:59]
  assign _T_132 = _T_125 ? _T_130 : _T_131; // @[LZD.scala 49:35]
  assign _T_134 = {_T_127,_T_129,_T_132}; // @[Cat.scala 29:58]
  assign _T_135 = _T_73[3]; // @[Shift.scala 12:21]
  assign _T_136 = _T_134[3]; // @[Shift.scala 12:21]
  assign _T_137 = _T_135 | _T_136; // @[LZD.scala 49:16]
  assign _T_138 = ~ _T_136; // @[LZD.scala 49:27]
  assign _T_139 = _T_135 | _T_138; // @[LZD.scala 49:25]
  assign _T_140 = _T_73[2:0]; // @[LZD.scala 49:47]
  assign _T_141 = _T_134[2:0]; // @[LZD.scala 49:59]
  assign _T_142 = _T_135 ? _T_140 : _T_141; // @[LZD.scala 49:35]
  assign _T_144 = {_T_137,_T_139,_T_142}; // @[Cat.scala 29:58]
  assign _T_145 = _T_11[15:0]; // @[LZD.scala 44:32]
  assign _T_146 = _T_145[15:8]; // @[LZD.scala 43:32]
  assign _T_147 = _T_146[7:4]; // @[LZD.scala 43:32]
  assign _T_148 = _T_147[3:2]; // @[LZD.scala 43:32]
  assign _T_149 = _T_148 != 2'h0; // @[LZD.scala 39:14]
  assign _T_150 = _T_148[1]; // @[LZD.scala 39:21]
  assign _T_151 = _T_148[0]; // @[LZD.scala 39:30]
  assign _T_152 = ~ _T_151; // @[LZD.scala 39:27]
  assign _T_153 = _T_150 | _T_152; // @[LZD.scala 39:25]
  assign _T_154 = {_T_149,_T_153}; // @[Cat.scala 29:58]
  assign _T_155 = _T_147[1:0]; // @[LZD.scala 44:32]
  assign _T_156 = _T_155 != 2'h0; // @[LZD.scala 39:14]
  assign _T_157 = _T_155[1]; // @[LZD.scala 39:21]
  assign _T_158 = _T_155[0]; // @[LZD.scala 39:30]
  assign _T_159 = ~ _T_158; // @[LZD.scala 39:27]
  assign _T_160 = _T_157 | _T_159; // @[LZD.scala 39:25]
  assign _T_161 = {_T_156,_T_160}; // @[Cat.scala 29:58]
  assign _T_162 = _T_154[1]; // @[Shift.scala 12:21]
  assign _T_163 = _T_161[1]; // @[Shift.scala 12:21]
  assign _T_164 = _T_162 | _T_163; // @[LZD.scala 49:16]
  assign _T_165 = ~ _T_163; // @[LZD.scala 49:27]
  assign _T_166 = _T_162 | _T_165; // @[LZD.scala 49:25]
  assign _T_167 = _T_154[0:0]; // @[LZD.scala 49:47]
  assign _T_168 = _T_161[0:0]; // @[LZD.scala 49:59]
  assign _T_169 = _T_162 ? _T_167 : _T_168; // @[LZD.scala 49:35]
  assign _T_171 = {_T_164,_T_166,_T_169}; // @[Cat.scala 29:58]
  assign _T_172 = _T_146[3:0]; // @[LZD.scala 44:32]
  assign _T_173 = _T_172[3:2]; // @[LZD.scala 43:32]
  assign _T_174 = _T_173 != 2'h0; // @[LZD.scala 39:14]
  assign _T_175 = _T_173[1]; // @[LZD.scala 39:21]
  assign _T_176 = _T_173[0]; // @[LZD.scala 39:30]
  assign _T_177 = ~ _T_176; // @[LZD.scala 39:27]
  assign _T_178 = _T_175 | _T_177; // @[LZD.scala 39:25]
  assign _T_179 = {_T_174,_T_178}; // @[Cat.scala 29:58]
  assign _T_180 = _T_172[1:0]; // @[LZD.scala 44:32]
  assign _T_181 = _T_180 != 2'h0; // @[LZD.scala 39:14]
  assign _T_182 = _T_180[1]; // @[LZD.scala 39:21]
  assign _T_183 = _T_180[0]; // @[LZD.scala 39:30]
  assign _T_184 = ~ _T_183; // @[LZD.scala 39:27]
  assign _T_185 = _T_182 | _T_184; // @[LZD.scala 39:25]
  assign _T_186 = {_T_181,_T_185}; // @[Cat.scala 29:58]
  assign _T_187 = _T_179[1]; // @[Shift.scala 12:21]
  assign _T_188 = _T_186[1]; // @[Shift.scala 12:21]
  assign _T_189 = _T_187 | _T_188; // @[LZD.scala 49:16]
  assign _T_190 = ~ _T_188; // @[LZD.scala 49:27]
  assign _T_191 = _T_187 | _T_190; // @[LZD.scala 49:25]
  assign _T_192 = _T_179[0:0]; // @[LZD.scala 49:47]
  assign _T_193 = _T_186[0:0]; // @[LZD.scala 49:59]
  assign _T_194 = _T_187 ? _T_192 : _T_193; // @[LZD.scala 49:35]
  assign _T_196 = {_T_189,_T_191,_T_194}; // @[Cat.scala 29:58]
  assign _T_197 = _T_171[2]; // @[Shift.scala 12:21]
  assign _T_198 = _T_196[2]; // @[Shift.scala 12:21]
  assign _T_199 = _T_197 | _T_198; // @[LZD.scala 49:16]
  assign _T_200 = ~ _T_198; // @[LZD.scala 49:27]
  assign _T_201 = _T_197 | _T_200; // @[LZD.scala 49:25]
  assign _T_202 = _T_171[1:0]; // @[LZD.scala 49:47]
  assign _T_203 = _T_196[1:0]; // @[LZD.scala 49:59]
  assign _T_204 = _T_197 ? _T_202 : _T_203; // @[LZD.scala 49:35]
  assign _T_206 = {_T_199,_T_201,_T_204}; // @[Cat.scala 29:58]
  assign _T_207 = _T_145[7:0]; // @[LZD.scala 44:32]
  assign _T_208 = _T_207[7:4]; // @[LZD.scala 43:32]
  assign _T_209 = _T_208[3:2]; // @[LZD.scala 43:32]
  assign _T_210 = _T_209 != 2'h0; // @[LZD.scala 39:14]
  assign _T_211 = _T_209[1]; // @[LZD.scala 39:21]
  assign _T_212 = _T_209[0]; // @[LZD.scala 39:30]
  assign _T_213 = ~ _T_212; // @[LZD.scala 39:27]
  assign _T_214 = _T_211 | _T_213; // @[LZD.scala 39:25]
  assign _T_215 = {_T_210,_T_214}; // @[Cat.scala 29:58]
  assign _T_216 = _T_208[1:0]; // @[LZD.scala 44:32]
  assign _T_217 = _T_216 != 2'h0; // @[LZD.scala 39:14]
  assign _T_218 = _T_216[1]; // @[LZD.scala 39:21]
  assign _T_219 = _T_216[0]; // @[LZD.scala 39:30]
  assign _T_220 = ~ _T_219; // @[LZD.scala 39:27]
  assign _T_221 = _T_218 | _T_220; // @[LZD.scala 39:25]
  assign _T_222 = {_T_217,_T_221}; // @[Cat.scala 29:58]
  assign _T_223 = _T_215[1]; // @[Shift.scala 12:21]
  assign _T_224 = _T_222[1]; // @[Shift.scala 12:21]
  assign _T_225 = _T_223 | _T_224; // @[LZD.scala 49:16]
  assign _T_226 = ~ _T_224; // @[LZD.scala 49:27]
  assign _T_227 = _T_223 | _T_226; // @[LZD.scala 49:25]
  assign _T_228 = _T_215[0:0]; // @[LZD.scala 49:47]
  assign _T_229 = _T_222[0:0]; // @[LZD.scala 49:59]
  assign _T_230 = _T_223 ? _T_228 : _T_229; // @[LZD.scala 49:35]
  assign _T_232 = {_T_225,_T_227,_T_230}; // @[Cat.scala 29:58]
  assign _T_233 = _T_207[3:0]; // @[LZD.scala 44:32]
  assign _T_234 = _T_233[3:2]; // @[LZD.scala 43:32]
  assign _T_235 = _T_234 != 2'h0; // @[LZD.scala 39:14]
  assign _T_236 = _T_234[1]; // @[LZD.scala 39:21]
  assign _T_237 = _T_234[0]; // @[LZD.scala 39:30]
  assign _T_238 = ~ _T_237; // @[LZD.scala 39:27]
  assign _T_239 = _T_236 | _T_238; // @[LZD.scala 39:25]
  assign _T_240 = {_T_235,_T_239}; // @[Cat.scala 29:58]
  assign _T_241 = _T_233[1:0]; // @[LZD.scala 44:32]
  assign _T_242 = _T_241 != 2'h0; // @[LZD.scala 39:14]
  assign _T_243 = _T_241[1]; // @[LZD.scala 39:21]
  assign _T_244 = _T_241[0]; // @[LZD.scala 39:30]
  assign _T_245 = ~ _T_244; // @[LZD.scala 39:27]
  assign _T_246 = _T_243 | _T_245; // @[LZD.scala 39:25]
  assign _T_247 = {_T_242,_T_246}; // @[Cat.scala 29:58]
  assign _T_248 = _T_240[1]; // @[Shift.scala 12:21]
  assign _T_249 = _T_247[1]; // @[Shift.scala 12:21]
  assign _T_250 = _T_248 | _T_249; // @[LZD.scala 49:16]
  assign _T_251 = ~ _T_249; // @[LZD.scala 49:27]
  assign _T_252 = _T_248 | _T_251; // @[LZD.scala 49:25]
  assign _T_253 = _T_240[0:0]; // @[LZD.scala 49:47]
  assign _T_254 = _T_247[0:0]; // @[LZD.scala 49:59]
  assign _T_255 = _T_248 ? _T_253 : _T_254; // @[LZD.scala 49:35]
  assign _T_257 = {_T_250,_T_252,_T_255}; // @[Cat.scala 29:58]
  assign _T_258 = _T_232[2]; // @[Shift.scala 12:21]
  assign _T_259 = _T_257[2]; // @[Shift.scala 12:21]
  assign _T_260 = _T_258 | _T_259; // @[LZD.scala 49:16]
  assign _T_261 = ~ _T_259; // @[LZD.scala 49:27]
  assign _T_262 = _T_258 | _T_261; // @[LZD.scala 49:25]
  assign _T_263 = _T_232[1:0]; // @[LZD.scala 49:47]
  assign _T_264 = _T_257[1:0]; // @[LZD.scala 49:59]
  assign _T_265 = _T_258 ? _T_263 : _T_264; // @[LZD.scala 49:35]
  assign _T_267 = {_T_260,_T_262,_T_265}; // @[Cat.scala 29:58]
  assign _T_268 = _T_206[3]; // @[Shift.scala 12:21]
  assign _T_269 = _T_267[3]; // @[Shift.scala 12:21]
  assign _T_270 = _T_268 | _T_269; // @[LZD.scala 49:16]
  assign _T_271 = ~ _T_269; // @[LZD.scala 49:27]
  assign _T_272 = _T_268 | _T_271; // @[LZD.scala 49:25]
  assign _T_273 = _T_206[2:0]; // @[LZD.scala 49:47]
  assign _T_274 = _T_267[2:0]; // @[LZD.scala 49:59]
  assign _T_275 = _T_268 ? _T_273 : _T_274; // @[LZD.scala 49:35]
  assign _T_277 = {_T_270,_T_272,_T_275}; // @[Cat.scala 29:58]
  assign _T_278 = _T_144[4]; // @[Shift.scala 12:21]
  assign _T_279 = _T_277[4]; // @[Shift.scala 12:21]
  assign _T_280 = _T_278 | _T_279; // @[LZD.scala 49:16]
  assign _T_281 = ~ _T_279; // @[LZD.scala 49:27]
  assign _T_282 = _T_278 | _T_281; // @[LZD.scala 49:25]
  assign _T_283 = _T_144[3:0]; // @[LZD.scala 49:47]
  assign _T_284 = _T_277[3:0]; // @[LZD.scala 49:59]
  assign _T_285 = _T_278 ? _T_283 : _T_284; // @[LZD.scala 49:35]
  assign _T_287 = {_T_280,_T_282,_T_285}; // @[Cat.scala 29:58]
  assign _T_288 = _T_10[31:0]; // @[LZD.scala 44:32]
  assign _T_289 = _T_288[31:16]; // @[LZD.scala 43:32]
  assign _T_290 = _T_289[15:8]; // @[LZD.scala 43:32]
  assign _T_291 = _T_290[7:4]; // @[LZD.scala 43:32]
  assign _T_292 = _T_291[3:2]; // @[LZD.scala 43:32]
  assign _T_293 = _T_292 != 2'h0; // @[LZD.scala 39:14]
  assign _T_294 = _T_292[1]; // @[LZD.scala 39:21]
  assign _T_295 = _T_292[0]; // @[LZD.scala 39:30]
  assign _T_296 = ~ _T_295; // @[LZD.scala 39:27]
  assign _T_297 = _T_294 | _T_296; // @[LZD.scala 39:25]
  assign _T_298 = {_T_293,_T_297}; // @[Cat.scala 29:58]
  assign _T_299 = _T_291[1:0]; // @[LZD.scala 44:32]
  assign _T_300 = _T_299 != 2'h0; // @[LZD.scala 39:14]
  assign _T_301 = _T_299[1]; // @[LZD.scala 39:21]
  assign _T_302 = _T_299[0]; // @[LZD.scala 39:30]
  assign _T_303 = ~ _T_302; // @[LZD.scala 39:27]
  assign _T_304 = _T_301 | _T_303; // @[LZD.scala 39:25]
  assign _T_305 = {_T_300,_T_304}; // @[Cat.scala 29:58]
  assign _T_306 = _T_298[1]; // @[Shift.scala 12:21]
  assign _T_307 = _T_305[1]; // @[Shift.scala 12:21]
  assign _T_308 = _T_306 | _T_307; // @[LZD.scala 49:16]
  assign _T_309 = ~ _T_307; // @[LZD.scala 49:27]
  assign _T_310 = _T_306 | _T_309; // @[LZD.scala 49:25]
  assign _T_311 = _T_298[0:0]; // @[LZD.scala 49:47]
  assign _T_312 = _T_305[0:0]; // @[LZD.scala 49:59]
  assign _T_313 = _T_306 ? _T_311 : _T_312; // @[LZD.scala 49:35]
  assign _T_315 = {_T_308,_T_310,_T_313}; // @[Cat.scala 29:58]
  assign _T_316 = _T_290[3:0]; // @[LZD.scala 44:32]
  assign _T_317 = _T_316[3:2]; // @[LZD.scala 43:32]
  assign _T_318 = _T_317 != 2'h0; // @[LZD.scala 39:14]
  assign _T_319 = _T_317[1]; // @[LZD.scala 39:21]
  assign _T_320 = _T_317[0]; // @[LZD.scala 39:30]
  assign _T_321 = ~ _T_320; // @[LZD.scala 39:27]
  assign _T_322 = _T_319 | _T_321; // @[LZD.scala 39:25]
  assign _T_323 = {_T_318,_T_322}; // @[Cat.scala 29:58]
  assign _T_324 = _T_316[1:0]; // @[LZD.scala 44:32]
  assign _T_325 = _T_324 != 2'h0; // @[LZD.scala 39:14]
  assign _T_326 = _T_324[1]; // @[LZD.scala 39:21]
  assign _T_327 = _T_324[0]; // @[LZD.scala 39:30]
  assign _T_328 = ~ _T_327; // @[LZD.scala 39:27]
  assign _T_329 = _T_326 | _T_328; // @[LZD.scala 39:25]
  assign _T_330 = {_T_325,_T_329}; // @[Cat.scala 29:58]
  assign _T_331 = _T_323[1]; // @[Shift.scala 12:21]
  assign _T_332 = _T_330[1]; // @[Shift.scala 12:21]
  assign _T_333 = _T_331 | _T_332; // @[LZD.scala 49:16]
  assign _T_334 = ~ _T_332; // @[LZD.scala 49:27]
  assign _T_335 = _T_331 | _T_334; // @[LZD.scala 49:25]
  assign _T_336 = _T_323[0:0]; // @[LZD.scala 49:47]
  assign _T_337 = _T_330[0:0]; // @[LZD.scala 49:59]
  assign _T_338 = _T_331 ? _T_336 : _T_337; // @[LZD.scala 49:35]
  assign _T_340 = {_T_333,_T_335,_T_338}; // @[Cat.scala 29:58]
  assign _T_341 = _T_315[2]; // @[Shift.scala 12:21]
  assign _T_342 = _T_340[2]; // @[Shift.scala 12:21]
  assign _T_343 = _T_341 | _T_342; // @[LZD.scala 49:16]
  assign _T_344 = ~ _T_342; // @[LZD.scala 49:27]
  assign _T_345 = _T_341 | _T_344; // @[LZD.scala 49:25]
  assign _T_346 = _T_315[1:0]; // @[LZD.scala 49:47]
  assign _T_347 = _T_340[1:0]; // @[LZD.scala 49:59]
  assign _T_348 = _T_341 ? _T_346 : _T_347; // @[LZD.scala 49:35]
  assign _T_350 = {_T_343,_T_345,_T_348}; // @[Cat.scala 29:58]
  assign _T_351 = _T_289[7:0]; // @[LZD.scala 44:32]
  assign _T_352 = _T_351[7:4]; // @[LZD.scala 43:32]
  assign _T_353 = _T_352[3:2]; // @[LZD.scala 43:32]
  assign _T_354 = _T_353 != 2'h0; // @[LZD.scala 39:14]
  assign _T_355 = _T_353[1]; // @[LZD.scala 39:21]
  assign _T_356 = _T_353[0]; // @[LZD.scala 39:30]
  assign _T_357 = ~ _T_356; // @[LZD.scala 39:27]
  assign _T_358 = _T_355 | _T_357; // @[LZD.scala 39:25]
  assign _T_359 = {_T_354,_T_358}; // @[Cat.scala 29:58]
  assign _T_360 = _T_352[1:0]; // @[LZD.scala 44:32]
  assign _T_361 = _T_360 != 2'h0; // @[LZD.scala 39:14]
  assign _T_362 = _T_360[1]; // @[LZD.scala 39:21]
  assign _T_363 = _T_360[0]; // @[LZD.scala 39:30]
  assign _T_364 = ~ _T_363; // @[LZD.scala 39:27]
  assign _T_365 = _T_362 | _T_364; // @[LZD.scala 39:25]
  assign _T_366 = {_T_361,_T_365}; // @[Cat.scala 29:58]
  assign _T_367 = _T_359[1]; // @[Shift.scala 12:21]
  assign _T_368 = _T_366[1]; // @[Shift.scala 12:21]
  assign _T_369 = _T_367 | _T_368; // @[LZD.scala 49:16]
  assign _T_370 = ~ _T_368; // @[LZD.scala 49:27]
  assign _T_371 = _T_367 | _T_370; // @[LZD.scala 49:25]
  assign _T_372 = _T_359[0:0]; // @[LZD.scala 49:47]
  assign _T_373 = _T_366[0:0]; // @[LZD.scala 49:59]
  assign _T_374 = _T_367 ? _T_372 : _T_373; // @[LZD.scala 49:35]
  assign _T_376 = {_T_369,_T_371,_T_374}; // @[Cat.scala 29:58]
  assign _T_377 = _T_351[3:0]; // @[LZD.scala 44:32]
  assign _T_378 = _T_377[3:2]; // @[LZD.scala 43:32]
  assign _T_379 = _T_378 != 2'h0; // @[LZD.scala 39:14]
  assign _T_380 = _T_378[1]; // @[LZD.scala 39:21]
  assign _T_381 = _T_378[0]; // @[LZD.scala 39:30]
  assign _T_382 = ~ _T_381; // @[LZD.scala 39:27]
  assign _T_383 = _T_380 | _T_382; // @[LZD.scala 39:25]
  assign _T_384 = {_T_379,_T_383}; // @[Cat.scala 29:58]
  assign _T_385 = _T_377[1:0]; // @[LZD.scala 44:32]
  assign _T_386 = _T_385 != 2'h0; // @[LZD.scala 39:14]
  assign _T_387 = _T_385[1]; // @[LZD.scala 39:21]
  assign _T_388 = _T_385[0]; // @[LZD.scala 39:30]
  assign _T_389 = ~ _T_388; // @[LZD.scala 39:27]
  assign _T_390 = _T_387 | _T_389; // @[LZD.scala 39:25]
  assign _T_391 = {_T_386,_T_390}; // @[Cat.scala 29:58]
  assign _T_392 = _T_384[1]; // @[Shift.scala 12:21]
  assign _T_393 = _T_391[1]; // @[Shift.scala 12:21]
  assign _T_394 = _T_392 | _T_393; // @[LZD.scala 49:16]
  assign _T_395 = ~ _T_393; // @[LZD.scala 49:27]
  assign _T_396 = _T_392 | _T_395; // @[LZD.scala 49:25]
  assign _T_397 = _T_384[0:0]; // @[LZD.scala 49:47]
  assign _T_398 = _T_391[0:0]; // @[LZD.scala 49:59]
  assign _T_399 = _T_392 ? _T_397 : _T_398; // @[LZD.scala 49:35]
  assign _T_401 = {_T_394,_T_396,_T_399}; // @[Cat.scala 29:58]
  assign _T_402 = _T_376[2]; // @[Shift.scala 12:21]
  assign _T_403 = _T_401[2]; // @[Shift.scala 12:21]
  assign _T_404 = _T_402 | _T_403; // @[LZD.scala 49:16]
  assign _T_405 = ~ _T_403; // @[LZD.scala 49:27]
  assign _T_406 = _T_402 | _T_405; // @[LZD.scala 49:25]
  assign _T_407 = _T_376[1:0]; // @[LZD.scala 49:47]
  assign _T_408 = _T_401[1:0]; // @[LZD.scala 49:59]
  assign _T_409 = _T_402 ? _T_407 : _T_408; // @[LZD.scala 49:35]
  assign _T_411 = {_T_404,_T_406,_T_409}; // @[Cat.scala 29:58]
  assign _T_412 = _T_350[3]; // @[Shift.scala 12:21]
  assign _T_413 = _T_411[3]; // @[Shift.scala 12:21]
  assign _T_414 = _T_412 | _T_413; // @[LZD.scala 49:16]
  assign _T_415 = ~ _T_413; // @[LZD.scala 49:27]
  assign _T_416 = _T_412 | _T_415; // @[LZD.scala 49:25]
  assign _T_417 = _T_350[2:0]; // @[LZD.scala 49:47]
  assign _T_418 = _T_411[2:0]; // @[LZD.scala 49:59]
  assign _T_419 = _T_412 ? _T_417 : _T_418; // @[LZD.scala 49:35]
  assign _T_421 = {_T_414,_T_416,_T_419}; // @[Cat.scala 29:58]
  assign _T_422 = _T_288[15:0]; // @[LZD.scala 44:32]
  assign _T_423 = _T_422[15:8]; // @[LZD.scala 43:32]
  assign _T_424 = _T_423[7:4]; // @[LZD.scala 43:32]
  assign _T_425 = _T_424[3:2]; // @[LZD.scala 43:32]
  assign _T_426 = _T_425 != 2'h0; // @[LZD.scala 39:14]
  assign _T_427 = _T_425[1]; // @[LZD.scala 39:21]
  assign _T_428 = _T_425[0]; // @[LZD.scala 39:30]
  assign _T_429 = ~ _T_428; // @[LZD.scala 39:27]
  assign _T_430 = _T_427 | _T_429; // @[LZD.scala 39:25]
  assign _T_431 = {_T_426,_T_430}; // @[Cat.scala 29:58]
  assign _T_432 = _T_424[1:0]; // @[LZD.scala 44:32]
  assign _T_433 = _T_432 != 2'h0; // @[LZD.scala 39:14]
  assign _T_434 = _T_432[1]; // @[LZD.scala 39:21]
  assign _T_435 = _T_432[0]; // @[LZD.scala 39:30]
  assign _T_436 = ~ _T_435; // @[LZD.scala 39:27]
  assign _T_437 = _T_434 | _T_436; // @[LZD.scala 39:25]
  assign _T_438 = {_T_433,_T_437}; // @[Cat.scala 29:58]
  assign _T_439 = _T_431[1]; // @[Shift.scala 12:21]
  assign _T_440 = _T_438[1]; // @[Shift.scala 12:21]
  assign _T_441 = _T_439 | _T_440; // @[LZD.scala 49:16]
  assign _T_442 = ~ _T_440; // @[LZD.scala 49:27]
  assign _T_443 = _T_439 | _T_442; // @[LZD.scala 49:25]
  assign _T_444 = _T_431[0:0]; // @[LZD.scala 49:47]
  assign _T_445 = _T_438[0:0]; // @[LZD.scala 49:59]
  assign _T_446 = _T_439 ? _T_444 : _T_445; // @[LZD.scala 49:35]
  assign _T_448 = {_T_441,_T_443,_T_446}; // @[Cat.scala 29:58]
  assign _T_449 = _T_423[3:0]; // @[LZD.scala 44:32]
  assign _T_450 = _T_449[3:2]; // @[LZD.scala 43:32]
  assign _T_451 = _T_450 != 2'h0; // @[LZD.scala 39:14]
  assign _T_452 = _T_450[1]; // @[LZD.scala 39:21]
  assign _T_453 = _T_450[0]; // @[LZD.scala 39:30]
  assign _T_454 = ~ _T_453; // @[LZD.scala 39:27]
  assign _T_455 = _T_452 | _T_454; // @[LZD.scala 39:25]
  assign _T_456 = {_T_451,_T_455}; // @[Cat.scala 29:58]
  assign _T_457 = _T_449[1:0]; // @[LZD.scala 44:32]
  assign _T_458 = _T_457 != 2'h0; // @[LZD.scala 39:14]
  assign _T_459 = _T_457[1]; // @[LZD.scala 39:21]
  assign _T_460 = _T_457[0]; // @[LZD.scala 39:30]
  assign _T_461 = ~ _T_460; // @[LZD.scala 39:27]
  assign _T_462 = _T_459 | _T_461; // @[LZD.scala 39:25]
  assign _T_463 = {_T_458,_T_462}; // @[Cat.scala 29:58]
  assign _T_464 = _T_456[1]; // @[Shift.scala 12:21]
  assign _T_465 = _T_463[1]; // @[Shift.scala 12:21]
  assign _T_466 = _T_464 | _T_465; // @[LZD.scala 49:16]
  assign _T_467 = ~ _T_465; // @[LZD.scala 49:27]
  assign _T_468 = _T_464 | _T_467; // @[LZD.scala 49:25]
  assign _T_469 = _T_456[0:0]; // @[LZD.scala 49:47]
  assign _T_470 = _T_463[0:0]; // @[LZD.scala 49:59]
  assign _T_471 = _T_464 ? _T_469 : _T_470; // @[LZD.scala 49:35]
  assign _T_473 = {_T_466,_T_468,_T_471}; // @[Cat.scala 29:58]
  assign _T_474 = _T_448[2]; // @[Shift.scala 12:21]
  assign _T_475 = _T_473[2]; // @[Shift.scala 12:21]
  assign _T_476 = _T_474 | _T_475; // @[LZD.scala 49:16]
  assign _T_477 = ~ _T_475; // @[LZD.scala 49:27]
  assign _T_478 = _T_474 | _T_477; // @[LZD.scala 49:25]
  assign _T_479 = _T_448[1:0]; // @[LZD.scala 49:47]
  assign _T_480 = _T_473[1:0]; // @[LZD.scala 49:59]
  assign _T_481 = _T_474 ? _T_479 : _T_480; // @[LZD.scala 49:35]
  assign _T_483 = {_T_476,_T_478,_T_481}; // @[Cat.scala 29:58]
  assign _T_484 = _T_422[7:0]; // @[LZD.scala 44:32]
  assign _T_485 = _T_484[7:4]; // @[LZD.scala 43:32]
  assign _T_486 = _T_485[3:2]; // @[LZD.scala 43:32]
  assign _T_487 = _T_486 != 2'h0; // @[LZD.scala 39:14]
  assign _T_488 = _T_486[1]; // @[LZD.scala 39:21]
  assign _T_489 = _T_486[0]; // @[LZD.scala 39:30]
  assign _T_490 = ~ _T_489; // @[LZD.scala 39:27]
  assign _T_491 = _T_488 | _T_490; // @[LZD.scala 39:25]
  assign _T_492 = {_T_487,_T_491}; // @[Cat.scala 29:58]
  assign _T_493 = _T_485[1:0]; // @[LZD.scala 44:32]
  assign _T_494 = _T_493 != 2'h0; // @[LZD.scala 39:14]
  assign _T_495 = _T_493[1]; // @[LZD.scala 39:21]
  assign _T_496 = _T_493[0]; // @[LZD.scala 39:30]
  assign _T_497 = ~ _T_496; // @[LZD.scala 39:27]
  assign _T_498 = _T_495 | _T_497; // @[LZD.scala 39:25]
  assign _T_499 = {_T_494,_T_498}; // @[Cat.scala 29:58]
  assign _T_500 = _T_492[1]; // @[Shift.scala 12:21]
  assign _T_501 = _T_499[1]; // @[Shift.scala 12:21]
  assign _T_502 = _T_500 | _T_501; // @[LZD.scala 49:16]
  assign _T_503 = ~ _T_501; // @[LZD.scala 49:27]
  assign _T_504 = _T_500 | _T_503; // @[LZD.scala 49:25]
  assign _T_505 = _T_492[0:0]; // @[LZD.scala 49:47]
  assign _T_506 = _T_499[0:0]; // @[LZD.scala 49:59]
  assign _T_507 = _T_500 ? _T_505 : _T_506; // @[LZD.scala 49:35]
  assign _T_509 = {_T_502,_T_504,_T_507}; // @[Cat.scala 29:58]
  assign _T_510 = _T_484[3:0]; // @[LZD.scala 44:32]
  assign _T_511 = _T_510[3:2]; // @[LZD.scala 43:32]
  assign _T_512 = _T_511 != 2'h0; // @[LZD.scala 39:14]
  assign _T_513 = _T_511[1]; // @[LZD.scala 39:21]
  assign _T_514 = _T_511[0]; // @[LZD.scala 39:30]
  assign _T_515 = ~ _T_514; // @[LZD.scala 39:27]
  assign _T_516 = _T_513 | _T_515; // @[LZD.scala 39:25]
  assign _T_517 = {_T_512,_T_516}; // @[Cat.scala 29:58]
  assign _T_518 = _T_510[1:0]; // @[LZD.scala 44:32]
  assign _T_519 = _T_518 != 2'h0; // @[LZD.scala 39:14]
  assign _T_520 = _T_518[1]; // @[LZD.scala 39:21]
  assign _T_521 = _T_518[0]; // @[LZD.scala 39:30]
  assign _T_522 = ~ _T_521; // @[LZD.scala 39:27]
  assign _T_523 = _T_520 | _T_522; // @[LZD.scala 39:25]
  assign _T_524 = {_T_519,_T_523}; // @[Cat.scala 29:58]
  assign _T_525 = _T_517[1]; // @[Shift.scala 12:21]
  assign _T_526 = _T_524[1]; // @[Shift.scala 12:21]
  assign _T_527 = _T_525 | _T_526; // @[LZD.scala 49:16]
  assign _T_528 = ~ _T_526; // @[LZD.scala 49:27]
  assign _T_529 = _T_525 | _T_528; // @[LZD.scala 49:25]
  assign _T_530 = _T_517[0:0]; // @[LZD.scala 49:47]
  assign _T_531 = _T_524[0:0]; // @[LZD.scala 49:59]
  assign _T_532 = _T_525 ? _T_530 : _T_531; // @[LZD.scala 49:35]
  assign _T_534 = {_T_527,_T_529,_T_532}; // @[Cat.scala 29:58]
  assign _T_535 = _T_509[2]; // @[Shift.scala 12:21]
  assign _T_536 = _T_534[2]; // @[Shift.scala 12:21]
  assign _T_537 = _T_535 | _T_536; // @[LZD.scala 49:16]
  assign _T_538 = ~ _T_536; // @[LZD.scala 49:27]
  assign _T_539 = _T_535 | _T_538; // @[LZD.scala 49:25]
  assign _T_540 = _T_509[1:0]; // @[LZD.scala 49:47]
  assign _T_541 = _T_534[1:0]; // @[LZD.scala 49:59]
  assign _T_542 = _T_535 ? _T_540 : _T_541; // @[LZD.scala 49:35]
  assign _T_544 = {_T_537,_T_539,_T_542}; // @[Cat.scala 29:58]
  assign _T_545 = _T_483[3]; // @[Shift.scala 12:21]
  assign _T_546 = _T_544[3]; // @[Shift.scala 12:21]
  assign _T_547 = _T_545 | _T_546; // @[LZD.scala 49:16]
  assign _T_548 = ~ _T_546; // @[LZD.scala 49:27]
  assign _T_549 = _T_545 | _T_548; // @[LZD.scala 49:25]
  assign _T_550 = _T_483[2:0]; // @[LZD.scala 49:47]
  assign _T_551 = _T_544[2:0]; // @[LZD.scala 49:59]
  assign _T_552 = _T_545 ? _T_550 : _T_551; // @[LZD.scala 49:35]
  assign _T_554 = {_T_547,_T_549,_T_552}; // @[Cat.scala 29:58]
  assign _T_555 = _T_421[4]; // @[Shift.scala 12:21]
  assign _T_556 = _T_554[4]; // @[Shift.scala 12:21]
  assign _T_557 = _T_555 | _T_556; // @[LZD.scala 49:16]
  assign _T_558 = ~ _T_556; // @[LZD.scala 49:27]
  assign _T_559 = _T_555 | _T_558; // @[LZD.scala 49:25]
  assign _T_560 = _T_421[3:0]; // @[LZD.scala 49:47]
  assign _T_561 = _T_554[3:0]; // @[LZD.scala 49:59]
  assign _T_562 = _T_555 ? _T_560 : _T_561; // @[LZD.scala 49:35]
  assign _T_564 = {_T_557,_T_559,_T_562}; // @[Cat.scala 29:58]
  assign _T_565 = _T_287[5]; // @[Shift.scala 12:21]
  assign _T_566 = _T_564[5]; // @[Shift.scala 12:21]
  assign _T_567 = _T_565 | _T_566; // @[LZD.scala 49:16]
  assign _T_568 = ~ _T_566; // @[LZD.scala 49:27]
  assign _T_569 = _T_565 | _T_568; // @[LZD.scala 49:25]
  assign _T_570 = _T_287[4:0]; // @[LZD.scala 49:47]
  assign _T_571 = _T_564[4:0]; // @[LZD.scala 49:59]
  assign _T_572 = _T_565 ? _T_570 : _T_571; // @[LZD.scala 49:35]
  assign _T_574 = {_T_567,_T_569,_T_572}; // @[Cat.scala 29:58]
  assign _T_575 = quireXOR[62:0]; // @[LZD.scala 44:32]
  assign _T_576 = _T_575[62:31]; // @[LZD.scala 43:32]
  assign _T_577 = _T_576[31:16]; // @[LZD.scala 43:32]
  assign _T_578 = _T_577[15:8]; // @[LZD.scala 43:32]
  assign _T_579 = _T_578[7:4]; // @[LZD.scala 43:32]
  assign _T_580 = _T_579[3:2]; // @[LZD.scala 43:32]
  assign _T_581 = _T_580 != 2'h0; // @[LZD.scala 39:14]
  assign _T_582 = _T_580[1]; // @[LZD.scala 39:21]
  assign _T_583 = _T_580[0]; // @[LZD.scala 39:30]
  assign _T_584 = ~ _T_583; // @[LZD.scala 39:27]
  assign _T_585 = _T_582 | _T_584; // @[LZD.scala 39:25]
  assign _T_586 = {_T_581,_T_585}; // @[Cat.scala 29:58]
  assign _T_587 = _T_579[1:0]; // @[LZD.scala 44:32]
  assign _T_588 = _T_587 != 2'h0; // @[LZD.scala 39:14]
  assign _T_589 = _T_587[1]; // @[LZD.scala 39:21]
  assign _T_590 = _T_587[0]; // @[LZD.scala 39:30]
  assign _T_591 = ~ _T_590; // @[LZD.scala 39:27]
  assign _T_592 = _T_589 | _T_591; // @[LZD.scala 39:25]
  assign _T_593 = {_T_588,_T_592}; // @[Cat.scala 29:58]
  assign _T_594 = _T_586[1]; // @[Shift.scala 12:21]
  assign _T_595 = _T_593[1]; // @[Shift.scala 12:21]
  assign _T_596 = _T_594 | _T_595; // @[LZD.scala 49:16]
  assign _T_597 = ~ _T_595; // @[LZD.scala 49:27]
  assign _T_598 = _T_594 | _T_597; // @[LZD.scala 49:25]
  assign _T_599 = _T_586[0:0]; // @[LZD.scala 49:47]
  assign _T_600 = _T_593[0:0]; // @[LZD.scala 49:59]
  assign _T_601 = _T_594 ? _T_599 : _T_600; // @[LZD.scala 49:35]
  assign _T_603 = {_T_596,_T_598,_T_601}; // @[Cat.scala 29:58]
  assign _T_604 = _T_578[3:0]; // @[LZD.scala 44:32]
  assign _T_605 = _T_604[3:2]; // @[LZD.scala 43:32]
  assign _T_606 = _T_605 != 2'h0; // @[LZD.scala 39:14]
  assign _T_607 = _T_605[1]; // @[LZD.scala 39:21]
  assign _T_608 = _T_605[0]; // @[LZD.scala 39:30]
  assign _T_609 = ~ _T_608; // @[LZD.scala 39:27]
  assign _T_610 = _T_607 | _T_609; // @[LZD.scala 39:25]
  assign _T_611 = {_T_606,_T_610}; // @[Cat.scala 29:58]
  assign _T_612 = _T_604[1:0]; // @[LZD.scala 44:32]
  assign _T_613 = _T_612 != 2'h0; // @[LZD.scala 39:14]
  assign _T_614 = _T_612[1]; // @[LZD.scala 39:21]
  assign _T_615 = _T_612[0]; // @[LZD.scala 39:30]
  assign _T_616 = ~ _T_615; // @[LZD.scala 39:27]
  assign _T_617 = _T_614 | _T_616; // @[LZD.scala 39:25]
  assign _T_618 = {_T_613,_T_617}; // @[Cat.scala 29:58]
  assign _T_619 = _T_611[1]; // @[Shift.scala 12:21]
  assign _T_620 = _T_618[1]; // @[Shift.scala 12:21]
  assign _T_621 = _T_619 | _T_620; // @[LZD.scala 49:16]
  assign _T_622 = ~ _T_620; // @[LZD.scala 49:27]
  assign _T_623 = _T_619 | _T_622; // @[LZD.scala 49:25]
  assign _T_624 = _T_611[0:0]; // @[LZD.scala 49:47]
  assign _T_625 = _T_618[0:0]; // @[LZD.scala 49:59]
  assign _T_626 = _T_619 ? _T_624 : _T_625; // @[LZD.scala 49:35]
  assign _T_628 = {_T_621,_T_623,_T_626}; // @[Cat.scala 29:58]
  assign _T_629 = _T_603[2]; // @[Shift.scala 12:21]
  assign _T_630 = _T_628[2]; // @[Shift.scala 12:21]
  assign _T_631 = _T_629 | _T_630; // @[LZD.scala 49:16]
  assign _T_632 = ~ _T_630; // @[LZD.scala 49:27]
  assign _T_633 = _T_629 | _T_632; // @[LZD.scala 49:25]
  assign _T_634 = _T_603[1:0]; // @[LZD.scala 49:47]
  assign _T_635 = _T_628[1:0]; // @[LZD.scala 49:59]
  assign _T_636 = _T_629 ? _T_634 : _T_635; // @[LZD.scala 49:35]
  assign _T_638 = {_T_631,_T_633,_T_636}; // @[Cat.scala 29:58]
  assign _T_639 = _T_577[7:0]; // @[LZD.scala 44:32]
  assign _T_640 = _T_639[7:4]; // @[LZD.scala 43:32]
  assign _T_641 = _T_640[3:2]; // @[LZD.scala 43:32]
  assign _T_642 = _T_641 != 2'h0; // @[LZD.scala 39:14]
  assign _T_643 = _T_641[1]; // @[LZD.scala 39:21]
  assign _T_644 = _T_641[0]; // @[LZD.scala 39:30]
  assign _T_645 = ~ _T_644; // @[LZD.scala 39:27]
  assign _T_646 = _T_643 | _T_645; // @[LZD.scala 39:25]
  assign _T_647 = {_T_642,_T_646}; // @[Cat.scala 29:58]
  assign _T_648 = _T_640[1:0]; // @[LZD.scala 44:32]
  assign _T_649 = _T_648 != 2'h0; // @[LZD.scala 39:14]
  assign _T_650 = _T_648[1]; // @[LZD.scala 39:21]
  assign _T_651 = _T_648[0]; // @[LZD.scala 39:30]
  assign _T_652 = ~ _T_651; // @[LZD.scala 39:27]
  assign _T_653 = _T_650 | _T_652; // @[LZD.scala 39:25]
  assign _T_654 = {_T_649,_T_653}; // @[Cat.scala 29:58]
  assign _T_655 = _T_647[1]; // @[Shift.scala 12:21]
  assign _T_656 = _T_654[1]; // @[Shift.scala 12:21]
  assign _T_657 = _T_655 | _T_656; // @[LZD.scala 49:16]
  assign _T_658 = ~ _T_656; // @[LZD.scala 49:27]
  assign _T_659 = _T_655 | _T_658; // @[LZD.scala 49:25]
  assign _T_660 = _T_647[0:0]; // @[LZD.scala 49:47]
  assign _T_661 = _T_654[0:0]; // @[LZD.scala 49:59]
  assign _T_662 = _T_655 ? _T_660 : _T_661; // @[LZD.scala 49:35]
  assign _T_664 = {_T_657,_T_659,_T_662}; // @[Cat.scala 29:58]
  assign _T_665 = _T_639[3:0]; // @[LZD.scala 44:32]
  assign _T_666 = _T_665[3:2]; // @[LZD.scala 43:32]
  assign _T_667 = _T_666 != 2'h0; // @[LZD.scala 39:14]
  assign _T_668 = _T_666[1]; // @[LZD.scala 39:21]
  assign _T_669 = _T_666[0]; // @[LZD.scala 39:30]
  assign _T_670 = ~ _T_669; // @[LZD.scala 39:27]
  assign _T_671 = _T_668 | _T_670; // @[LZD.scala 39:25]
  assign _T_672 = {_T_667,_T_671}; // @[Cat.scala 29:58]
  assign _T_673 = _T_665[1:0]; // @[LZD.scala 44:32]
  assign _T_674 = _T_673 != 2'h0; // @[LZD.scala 39:14]
  assign _T_675 = _T_673[1]; // @[LZD.scala 39:21]
  assign _T_676 = _T_673[0]; // @[LZD.scala 39:30]
  assign _T_677 = ~ _T_676; // @[LZD.scala 39:27]
  assign _T_678 = _T_675 | _T_677; // @[LZD.scala 39:25]
  assign _T_679 = {_T_674,_T_678}; // @[Cat.scala 29:58]
  assign _T_680 = _T_672[1]; // @[Shift.scala 12:21]
  assign _T_681 = _T_679[1]; // @[Shift.scala 12:21]
  assign _T_682 = _T_680 | _T_681; // @[LZD.scala 49:16]
  assign _T_683 = ~ _T_681; // @[LZD.scala 49:27]
  assign _T_684 = _T_680 | _T_683; // @[LZD.scala 49:25]
  assign _T_685 = _T_672[0:0]; // @[LZD.scala 49:47]
  assign _T_686 = _T_679[0:0]; // @[LZD.scala 49:59]
  assign _T_687 = _T_680 ? _T_685 : _T_686; // @[LZD.scala 49:35]
  assign _T_689 = {_T_682,_T_684,_T_687}; // @[Cat.scala 29:58]
  assign _T_690 = _T_664[2]; // @[Shift.scala 12:21]
  assign _T_691 = _T_689[2]; // @[Shift.scala 12:21]
  assign _T_692 = _T_690 | _T_691; // @[LZD.scala 49:16]
  assign _T_693 = ~ _T_691; // @[LZD.scala 49:27]
  assign _T_694 = _T_690 | _T_693; // @[LZD.scala 49:25]
  assign _T_695 = _T_664[1:0]; // @[LZD.scala 49:47]
  assign _T_696 = _T_689[1:0]; // @[LZD.scala 49:59]
  assign _T_697 = _T_690 ? _T_695 : _T_696; // @[LZD.scala 49:35]
  assign _T_699 = {_T_692,_T_694,_T_697}; // @[Cat.scala 29:58]
  assign _T_700 = _T_638[3]; // @[Shift.scala 12:21]
  assign _T_701 = _T_699[3]; // @[Shift.scala 12:21]
  assign _T_702 = _T_700 | _T_701; // @[LZD.scala 49:16]
  assign _T_703 = ~ _T_701; // @[LZD.scala 49:27]
  assign _T_704 = _T_700 | _T_703; // @[LZD.scala 49:25]
  assign _T_705 = _T_638[2:0]; // @[LZD.scala 49:47]
  assign _T_706 = _T_699[2:0]; // @[LZD.scala 49:59]
  assign _T_707 = _T_700 ? _T_705 : _T_706; // @[LZD.scala 49:35]
  assign _T_709 = {_T_702,_T_704,_T_707}; // @[Cat.scala 29:58]
  assign _T_710 = _T_576[15:0]; // @[LZD.scala 44:32]
  assign _T_711 = _T_710[15:8]; // @[LZD.scala 43:32]
  assign _T_712 = _T_711[7:4]; // @[LZD.scala 43:32]
  assign _T_713 = _T_712[3:2]; // @[LZD.scala 43:32]
  assign _T_714 = _T_713 != 2'h0; // @[LZD.scala 39:14]
  assign _T_715 = _T_713[1]; // @[LZD.scala 39:21]
  assign _T_716 = _T_713[0]; // @[LZD.scala 39:30]
  assign _T_717 = ~ _T_716; // @[LZD.scala 39:27]
  assign _T_718 = _T_715 | _T_717; // @[LZD.scala 39:25]
  assign _T_719 = {_T_714,_T_718}; // @[Cat.scala 29:58]
  assign _T_720 = _T_712[1:0]; // @[LZD.scala 44:32]
  assign _T_721 = _T_720 != 2'h0; // @[LZD.scala 39:14]
  assign _T_722 = _T_720[1]; // @[LZD.scala 39:21]
  assign _T_723 = _T_720[0]; // @[LZD.scala 39:30]
  assign _T_724 = ~ _T_723; // @[LZD.scala 39:27]
  assign _T_725 = _T_722 | _T_724; // @[LZD.scala 39:25]
  assign _T_726 = {_T_721,_T_725}; // @[Cat.scala 29:58]
  assign _T_727 = _T_719[1]; // @[Shift.scala 12:21]
  assign _T_728 = _T_726[1]; // @[Shift.scala 12:21]
  assign _T_729 = _T_727 | _T_728; // @[LZD.scala 49:16]
  assign _T_730 = ~ _T_728; // @[LZD.scala 49:27]
  assign _T_731 = _T_727 | _T_730; // @[LZD.scala 49:25]
  assign _T_732 = _T_719[0:0]; // @[LZD.scala 49:47]
  assign _T_733 = _T_726[0:0]; // @[LZD.scala 49:59]
  assign _T_734 = _T_727 ? _T_732 : _T_733; // @[LZD.scala 49:35]
  assign _T_736 = {_T_729,_T_731,_T_734}; // @[Cat.scala 29:58]
  assign _T_737 = _T_711[3:0]; // @[LZD.scala 44:32]
  assign _T_738 = _T_737[3:2]; // @[LZD.scala 43:32]
  assign _T_739 = _T_738 != 2'h0; // @[LZD.scala 39:14]
  assign _T_740 = _T_738[1]; // @[LZD.scala 39:21]
  assign _T_741 = _T_738[0]; // @[LZD.scala 39:30]
  assign _T_742 = ~ _T_741; // @[LZD.scala 39:27]
  assign _T_743 = _T_740 | _T_742; // @[LZD.scala 39:25]
  assign _T_744 = {_T_739,_T_743}; // @[Cat.scala 29:58]
  assign _T_745 = _T_737[1:0]; // @[LZD.scala 44:32]
  assign _T_746 = _T_745 != 2'h0; // @[LZD.scala 39:14]
  assign _T_747 = _T_745[1]; // @[LZD.scala 39:21]
  assign _T_748 = _T_745[0]; // @[LZD.scala 39:30]
  assign _T_749 = ~ _T_748; // @[LZD.scala 39:27]
  assign _T_750 = _T_747 | _T_749; // @[LZD.scala 39:25]
  assign _T_751 = {_T_746,_T_750}; // @[Cat.scala 29:58]
  assign _T_752 = _T_744[1]; // @[Shift.scala 12:21]
  assign _T_753 = _T_751[1]; // @[Shift.scala 12:21]
  assign _T_754 = _T_752 | _T_753; // @[LZD.scala 49:16]
  assign _T_755 = ~ _T_753; // @[LZD.scala 49:27]
  assign _T_756 = _T_752 | _T_755; // @[LZD.scala 49:25]
  assign _T_757 = _T_744[0:0]; // @[LZD.scala 49:47]
  assign _T_758 = _T_751[0:0]; // @[LZD.scala 49:59]
  assign _T_759 = _T_752 ? _T_757 : _T_758; // @[LZD.scala 49:35]
  assign _T_761 = {_T_754,_T_756,_T_759}; // @[Cat.scala 29:58]
  assign _T_762 = _T_736[2]; // @[Shift.scala 12:21]
  assign _T_763 = _T_761[2]; // @[Shift.scala 12:21]
  assign _T_764 = _T_762 | _T_763; // @[LZD.scala 49:16]
  assign _T_765 = ~ _T_763; // @[LZD.scala 49:27]
  assign _T_766 = _T_762 | _T_765; // @[LZD.scala 49:25]
  assign _T_767 = _T_736[1:0]; // @[LZD.scala 49:47]
  assign _T_768 = _T_761[1:0]; // @[LZD.scala 49:59]
  assign _T_769 = _T_762 ? _T_767 : _T_768; // @[LZD.scala 49:35]
  assign _T_771 = {_T_764,_T_766,_T_769}; // @[Cat.scala 29:58]
  assign _T_772 = _T_710[7:0]; // @[LZD.scala 44:32]
  assign _T_773 = _T_772[7:4]; // @[LZD.scala 43:32]
  assign _T_774 = _T_773[3:2]; // @[LZD.scala 43:32]
  assign _T_775 = _T_774 != 2'h0; // @[LZD.scala 39:14]
  assign _T_776 = _T_774[1]; // @[LZD.scala 39:21]
  assign _T_777 = _T_774[0]; // @[LZD.scala 39:30]
  assign _T_778 = ~ _T_777; // @[LZD.scala 39:27]
  assign _T_779 = _T_776 | _T_778; // @[LZD.scala 39:25]
  assign _T_780 = {_T_775,_T_779}; // @[Cat.scala 29:58]
  assign _T_781 = _T_773[1:0]; // @[LZD.scala 44:32]
  assign _T_782 = _T_781 != 2'h0; // @[LZD.scala 39:14]
  assign _T_783 = _T_781[1]; // @[LZD.scala 39:21]
  assign _T_784 = _T_781[0]; // @[LZD.scala 39:30]
  assign _T_785 = ~ _T_784; // @[LZD.scala 39:27]
  assign _T_786 = _T_783 | _T_785; // @[LZD.scala 39:25]
  assign _T_787 = {_T_782,_T_786}; // @[Cat.scala 29:58]
  assign _T_788 = _T_780[1]; // @[Shift.scala 12:21]
  assign _T_789 = _T_787[1]; // @[Shift.scala 12:21]
  assign _T_790 = _T_788 | _T_789; // @[LZD.scala 49:16]
  assign _T_791 = ~ _T_789; // @[LZD.scala 49:27]
  assign _T_792 = _T_788 | _T_791; // @[LZD.scala 49:25]
  assign _T_793 = _T_780[0:0]; // @[LZD.scala 49:47]
  assign _T_794 = _T_787[0:0]; // @[LZD.scala 49:59]
  assign _T_795 = _T_788 ? _T_793 : _T_794; // @[LZD.scala 49:35]
  assign _T_797 = {_T_790,_T_792,_T_795}; // @[Cat.scala 29:58]
  assign _T_798 = _T_772[3:0]; // @[LZD.scala 44:32]
  assign _T_799 = _T_798[3:2]; // @[LZD.scala 43:32]
  assign _T_800 = _T_799 != 2'h0; // @[LZD.scala 39:14]
  assign _T_801 = _T_799[1]; // @[LZD.scala 39:21]
  assign _T_802 = _T_799[0]; // @[LZD.scala 39:30]
  assign _T_803 = ~ _T_802; // @[LZD.scala 39:27]
  assign _T_804 = _T_801 | _T_803; // @[LZD.scala 39:25]
  assign _T_805 = {_T_800,_T_804}; // @[Cat.scala 29:58]
  assign _T_806 = _T_798[1:0]; // @[LZD.scala 44:32]
  assign _T_807 = _T_806 != 2'h0; // @[LZD.scala 39:14]
  assign _T_808 = _T_806[1]; // @[LZD.scala 39:21]
  assign _T_809 = _T_806[0]; // @[LZD.scala 39:30]
  assign _T_810 = ~ _T_809; // @[LZD.scala 39:27]
  assign _T_811 = _T_808 | _T_810; // @[LZD.scala 39:25]
  assign _T_812 = {_T_807,_T_811}; // @[Cat.scala 29:58]
  assign _T_813 = _T_805[1]; // @[Shift.scala 12:21]
  assign _T_814 = _T_812[1]; // @[Shift.scala 12:21]
  assign _T_815 = _T_813 | _T_814; // @[LZD.scala 49:16]
  assign _T_816 = ~ _T_814; // @[LZD.scala 49:27]
  assign _T_817 = _T_813 | _T_816; // @[LZD.scala 49:25]
  assign _T_818 = _T_805[0:0]; // @[LZD.scala 49:47]
  assign _T_819 = _T_812[0:0]; // @[LZD.scala 49:59]
  assign _T_820 = _T_813 ? _T_818 : _T_819; // @[LZD.scala 49:35]
  assign _T_822 = {_T_815,_T_817,_T_820}; // @[Cat.scala 29:58]
  assign _T_823 = _T_797[2]; // @[Shift.scala 12:21]
  assign _T_824 = _T_822[2]; // @[Shift.scala 12:21]
  assign _T_825 = _T_823 | _T_824; // @[LZD.scala 49:16]
  assign _T_826 = ~ _T_824; // @[LZD.scala 49:27]
  assign _T_827 = _T_823 | _T_826; // @[LZD.scala 49:25]
  assign _T_828 = _T_797[1:0]; // @[LZD.scala 49:47]
  assign _T_829 = _T_822[1:0]; // @[LZD.scala 49:59]
  assign _T_830 = _T_823 ? _T_828 : _T_829; // @[LZD.scala 49:35]
  assign _T_832 = {_T_825,_T_827,_T_830}; // @[Cat.scala 29:58]
  assign _T_833 = _T_771[3]; // @[Shift.scala 12:21]
  assign _T_834 = _T_832[3]; // @[Shift.scala 12:21]
  assign _T_835 = _T_833 | _T_834; // @[LZD.scala 49:16]
  assign _T_836 = ~ _T_834; // @[LZD.scala 49:27]
  assign _T_837 = _T_833 | _T_836; // @[LZD.scala 49:25]
  assign _T_838 = _T_771[2:0]; // @[LZD.scala 49:47]
  assign _T_839 = _T_832[2:0]; // @[LZD.scala 49:59]
  assign _T_840 = _T_833 ? _T_838 : _T_839; // @[LZD.scala 49:35]
  assign _T_842 = {_T_835,_T_837,_T_840}; // @[Cat.scala 29:58]
  assign _T_843 = _T_709[4]; // @[Shift.scala 12:21]
  assign _T_844 = _T_842[4]; // @[Shift.scala 12:21]
  assign _T_845 = _T_843 | _T_844; // @[LZD.scala 49:16]
  assign _T_846 = ~ _T_844; // @[LZD.scala 49:27]
  assign _T_847 = _T_843 | _T_846; // @[LZD.scala 49:25]
  assign _T_848 = _T_709[3:0]; // @[LZD.scala 49:47]
  assign _T_849 = _T_842[3:0]; // @[LZD.scala 49:59]
  assign _T_850 = _T_843 ? _T_848 : _T_849; // @[LZD.scala 49:35]
  assign _T_852 = {_T_845,_T_847,_T_850}; // @[Cat.scala 29:58]
  assign _T_853 = _T_575[30:0]; // @[LZD.scala 44:32]
  assign _T_854 = _T_853[30:15]; // @[LZD.scala 43:32]
  assign _T_855 = _T_854[15:8]; // @[LZD.scala 43:32]
  assign _T_856 = _T_855[7:4]; // @[LZD.scala 43:32]
  assign _T_857 = _T_856[3:2]; // @[LZD.scala 43:32]
  assign _T_858 = _T_857 != 2'h0; // @[LZD.scala 39:14]
  assign _T_859 = _T_857[1]; // @[LZD.scala 39:21]
  assign _T_860 = _T_857[0]; // @[LZD.scala 39:30]
  assign _T_861 = ~ _T_860; // @[LZD.scala 39:27]
  assign _T_862 = _T_859 | _T_861; // @[LZD.scala 39:25]
  assign _T_863 = {_T_858,_T_862}; // @[Cat.scala 29:58]
  assign _T_864 = _T_856[1:0]; // @[LZD.scala 44:32]
  assign _T_865 = _T_864 != 2'h0; // @[LZD.scala 39:14]
  assign _T_866 = _T_864[1]; // @[LZD.scala 39:21]
  assign _T_867 = _T_864[0]; // @[LZD.scala 39:30]
  assign _T_868 = ~ _T_867; // @[LZD.scala 39:27]
  assign _T_869 = _T_866 | _T_868; // @[LZD.scala 39:25]
  assign _T_870 = {_T_865,_T_869}; // @[Cat.scala 29:58]
  assign _T_871 = _T_863[1]; // @[Shift.scala 12:21]
  assign _T_872 = _T_870[1]; // @[Shift.scala 12:21]
  assign _T_873 = _T_871 | _T_872; // @[LZD.scala 49:16]
  assign _T_874 = ~ _T_872; // @[LZD.scala 49:27]
  assign _T_875 = _T_871 | _T_874; // @[LZD.scala 49:25]
  assign _T_876 = _T_863[0:0]; // @[LZD.scala 49:47]
  assign _T_877 = _T_870[0:0]; // @[LZD.scala 49:59]
  assign _T_878 = _T_871 ? _T_876 : _T_877; // @[LZD.scala 49:35]
  assign _T_880 = {_T_873,_T_875,_T_878}; // @[Cat.scala 29:58]
  assign _T_881 = _T_855[3:0]; // @[LZD.scala 44:32]
  assign _T_882 = _T_881[3:2]; // @[LZD.scala 43:32]
  assign _T_883 = _T_882 != 2'h0; // @[LZD.scala 39:14]
  assign _T_884 = _T_882[1]; // @[LZD.scala 39:21]
  assign _T_885 = _T_882[0]; // @[LZD.scala 39:30]
  assign _T_886 = ~ _T_885; // @[LZD.scala 39:27]
  assign _T_887 = _T_884 | _T_886; // @[LZD.scala 39:25]
  assign _T_888 = {_T_883,_T_887}; // @[Cat.scala 29:58]
  assign _T_889 = _T_881[1:0]; // @[LZD.scala 44:32]
  assign _T_890 = _T_889 != 2'h0; // @[LZD.scala 39:14]
  assign _T_891 = _T_889[1]; // @[LZD.scala 39:21]
  assign _T_892 = _T_889[0]; // @[LZD.scala 39:30]
  assign _T_893 = ~ _T_892; // @[LZD.scala 39:27]
  assign _T_894 = _T_891 | _T_893; // @[LZD.scala 39:25]
  assign _T_895 = {_T_890,_T_894}; // @[Cat.scala 29:58]
  assign _T_896 = _T_888[1]; // @[Shift.scala 12:21]
  assign _T_897 = _T_895[1]; // @[Shift.scala 12:21]
  assign _T_898 = _T_896 | _T_897; // @[LZD.scala 49:16]
  assign _T_899 = ~ _T_897; // @[LZD.scala 49:27]
  assign _T_900 = _T_896 | _T_899; // @[LZD.scala 49:25]
  assign _T_901 = _T_888[0:0]; // @[LZD.scala 49:47]
  assign _T_902 = _T_895[0:0]; // @[LZD.scala 49:59]
  assign _T_903 = _T_896 ? _T_901 : _T_902; // @[LZD.scala 49:35]
  assign _T_905 = {_T_898,_T_900,_T_903}; // @[Cat.scala 29:58]
  assign _T_906 = _T_880[2]; // @[Shift.scala 12:21]
  assign _T_907 = _T_905[2]; // @[Shift.scala 12:21]
  assign _T_908 = _T_906 | _T_907; // @[LZD.scala 49:16]
  assign _T_909 = ~ _T_907; // @[LZD.scala 49:27]
  assign _T_910 = _T_906 | _T_909; // @[LZD.scala 49:25]
  assign _T_911 = _T_880[1:0]; // @[LZD.scala 49:47]
  assign _T_912 = _T_905[1:0]; // @[LZD.scala 49:59]
  assign _T_913 = _T_906 ? _T_911 : _T_912; // @[LZD.scala 49:35]
  assign _T_915 = {_T_908,_T_910,_T_913}; // @[Cat.scala 29:58]
  assign _T_916 = _T_854[7:0]; // @[LZD.scala 44:32]
  assign _T_917 = _T_916[7:4]; // @[LZD.scala 43:32]
  assign _T_918 = _T_917[3:2]; // @[LZD.scala 43:32]
  assign _T_919 = _T_918 != 2'h0; // @[LZD.scala 39:14]
  assign _T_920 = _T_918[1]; // @[LZD.scala 39:21]
  assign _T_921 = _T_918[0]; // @[LZD.scala 39:30]
  assign _T_922 = ~ _T_921; // @[LZD.scala 39:27]
  assign _T_923 = _T_920 | _T_922; // @[LZD.scala 39:25]
  assign _T_924 = {_T_919,_T_923}; // @[Cat.scala 29:58]
  assign _T_925 = _T_917[1:0]; // @[LZD.scala 44:32]
  assign _T_926 = _T_925 != 2'h0; // @[LZD.scala 39:14]
  assign _T_927 = _T_925[1]; // @[LZD.scala 39:21]
  assign _T_928 = _T_925[0]; // @[LZD.scala 39:30]
  assign _T_929 = ~ _T_928; // @[LZD.scala 39:27]
  assign _T_930 = _T_927 | _T_929; // @[LZD.scala 39:25]
  assign _T_931 = {_T_926,_T_930}; // @[Cat.scala 29:58]
  assign _T_932 = _T_924[1]; // @[Shift.scala 12:21]
  assign _T_933 = _T_931[1]; // @[Shift.scala 12:21]
  assign _T_934 = _T_932 | _T_933; // @[LZD.scala 49:16]
  assign _T_935 = ~ _T_933; // @[LZD.scala 49:27]
  assign _T_936 = _T_932 | _T_935; // @[LZD.scala 49:25]
  assign _T_937 = _T_924[0:0]; // @[LZD.scala 49:47]
  assign _T_938 = _T_931[0:0]; // @[LZD.scala 49:59]
  assign _T_939 = _T_932 ? _T_937 : _T_938; // @[LZD.scala 49:35]
  assign _T_941 = {_T_934,_T_936,_T_939}; // @[Cat.scala 29:58]
  assign _T_942 = _T_916[3:0]; // @[LZD.scala 44:32]
  assign _T_943 = _T_942[3:2]; // @[LZD.scala 43:32]
  assign _T_944 = _T_943 != 2'h0; // @[LZD.scala 39:14]
  assign _T_945 = _T_943[1]; // @[LZD.scala 39:21]
  assign _T_946 = _T_943[0]; // @[LZD.scala 39:30]
  assign _T_947 = ~ _T_946; // @[LZD.scala 39:27]
  assign _T_948 = _T_945 | _T_947; // @[LZD.scala 39:25]
  assign _T_949 = {_T_944,_T_948}; // @[Cat.scala 29:58]
  assign _T_950 = _T_942[1:0]; // @[LZD.scala 44:32]
  assign _T_951 = _T_950 != 2'h0; // @[LZD.scala 39:14]
  assign _T_952 = _T_950[1]; // @[LZD.scala 39:21]
  assign _T_953 = _T_950[0]; // @[LZD.scala 39:30]
  assign _T_954 = ~ _T_953; // @[LZD.scala 39:27]
  assign _T_955 = _T_952 | _T_954; // @[LZD.scala 39:25]
  assign _T_956 = {_T_951,_T_955}; // @[Cat.scala 29:58]
  assign _T_957 = _T_949[1]; // @[Shift.scala 12:21]
  assign _T_958 = _T_956[1]; // @[Shift.scala 12:21]
  assign _T_959 = _T_957 | _T_958; // @[LZD.scala 49:16]
  assign _T_960 = ~ _T_958; // @[LZD.scala 49:27]
  assign _T_961 = _T_957 | _T_960; // @[LZD.scala 49:25]
  assign _T_962 = _T_949[0:0]; // @[LZD.scala 49:47]
  assign _T_963 = _T_956[0:0]; // @[LZD.scala 49:59]
  assign _T_964 = _T_957 ? _T_962 : _T_963; // @[LZD.scala 49:35]
  assign _T_966 = {_T_959,_T_961,_T_964}; // @[Cat.scala 29:58]
  assign _T_967 = _T_941[2]; // @[Shift.scala 12:21]
  assign _T_968 = _T_966[2]; // @[Shift.scala 12:21]
  assign _T_969 = _T_967 | _T_968; // @[LZD.scala 49:16]
  assign _T_970 = ~ _T_968; // @[LZD.scala 49:27]
  assign _T_971 = _T_967 | _T_970; // @[LZD.scala 49:25]
  assign _T_972 = _T_941[1:0]; // @[LZD.scala 49:47]
  assign _T_973 = _T_966[1:0]; // @[LZD.scala 49:59]
  assign _T_974 = _T_967 ? _T_972 : _T_973; // @[LZD.scala 49:35]
  assign _T_976 = {_T_969,_T_971,_T_974}; // @[Cat.scala 29:58]
  assign _T_977 = _T_915[3]; // @[Shift.scala 12:21]
  assign _T_978 = _T_976[3]; // @[Shift.scala 12:21]
  assign _T_979 = _T_977 | _T_978; // @[LZD.scala 49:16]
  assign _T_980 = ~ _T_978; // @[LZD.scala 49:27]
  assign _T_981 = _T_977 | _T_980; // @[LZD.scala 49:25]
  assign _T_982 = _T_915[2:0]; // @[LZD.scala 49:47]
  assign _T_983 = _T_976[2:0]; // @[LZD.scala 49:59]
  assign _T_984 = _T_977 ? _T_982 : _T_983; // @[LZD.scala 49:35]
  assign _T_986 = {_T_979,_T_981,_T_984}; // @[Cat.scala 29:58]
  assign _T_987 = _T_853[14:0]; // @[LZD.scala 44:32]
  assign _T_988 = _T_987[14:7]; // @[LZD.scala 43:32]
  assign _T_989 = _T_988[7:4]; // @[LZD.scala 43:32]
  assign _T_990 = _T_989[3:2]; // @[LZD.scala 43:32]
  assign _T_991 = _T_990 != 2'h0; // @[LZD.scala 39:14]
  assign _T_992 = _T_990[1]; // @[LZD.scala 39:21]
  assign _T_993 = _T_990[0]; // @[LZD.scala 39:30]
  assign _T_994 = ~ _T_993; // @[LZD.scala 39:27]
  assign _T_995 = _T_992 | _T_994; // @[LZD.scala 39:25]
  assign _T_996 = {_T_991,_T_995}; // @[Cat.scala 29:58]
  assign _T_997 = _T_989[1:0]; // @[LZD.scala 44:32]
  assign _T_998 = _T_997 != 2'h0; // @[LZD.scala 39:14]
  assign _T_999 = _T_997[1]; // @[LZD.scala 39:21]
  assign _T_1000 = _T_997[0]; // @[LZD.scala 39:30]
  assign _T_1001 = ~ _T_1000; // @[LZD.scala 39:27]
  assign _T_1002 = _T_999 | _T_1001; // @[LZD.scala 39:25]
  assign _T_1003 = {_T_998,_T_1002}; // @[Cat.scala 29:58]
  assign _T_1004 = _T_996[1]; // @[Shift.scala 12:21]
  assign _T_1005 = _T_1003[1]; // @[Shift.scala 12:21]
  assign _T_1006 = _T_1004 | _T_1005; // @[LZD.scala 49:16]
  assign _T_1007 = ~ _T_1005; // @[LZD.scala 49:27]
  assign _T_1008 = _T_1004 | _T_1007; // @[LZD.scala 49:25]
  assign _T_1009 = _T_996[0:0]; // @[LZD.scala 49:47]
  assign _T_1010 = _T_1003[0:0]; // @[LZD.scala 49:59]
  assign _T_1011 = _T_1004 ? _T_1009 : _T_1010; // @[LZD.scala 49:35]
  assign _T_1013 = {_T_1006,_T_1008,_T_1011}; // @[Cat.scala 29:58]
  assign _T_1014 = _T_988[3:0]; // @[LZD.scala 44:32]
  assign _T_1015 = _T_1014[3:2]; // @[LZD.scala 43:32]
  assign _T_1016 = _T_1015 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1017 = _T_1015[1]; // @[LZD.scala 39:21]
  assign _T_1018 = _T_1015[0]; // @[LZD.scala 39:30]
  assign _T_1019 = ~ _T_1018; // @[LZD.scala 39:27]
  assign _T_1020 = _T_1017 | _T_1019; // @[LZD.scala 39:25]
  assign _T_1021 = {_T_1016,_T_1020}; // @[Cat.scala 29:58]
  assign _T_1022 = _T_1014[1:0]; // @[LZD.scala 44:32]
  assign _T_1023 = _T_1022 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1024 = _T_1022[1]; // @[LZD.scala 39:21]
  assign _T_1025 = _T_1022[0]; // @[LZD.scala 39:30]
  assign _T_1026 = ~ _T_1025; // @[LZD.scala 39:27]
  assign _T_1027 = _T_1024 | _T_1026; // @[LZD.scala 39:25]
  assign _T_1028 = {_T_1023,_T_1027}; // @[Cat.scala 29:58]
  assign _T_1029 = _T_1021[1]; // @[Shift.scala 12:21]
  assign _T_1030 = _T_1028[1]; // @[Shift.scala 12:21]
  assign _T_1031 = _T_1029 | _T_1030; // @[LZD.scala 49:16]
  assign _T_1032 = ~ _T_1030; // @[LZD.scala 49:27]
  assign _T_1033 = _T_1029 | _T_1032; // @[LZD.scala 49:25]
  assign _T_1034 = _T_1021[0:0]; // @[LZD.scala 49:47]
  assign _T_1035 = _T_1028[0:0]; // @[LZD.scala 49:59]
  assign _T_1036 = _T_1029 ? _T_1034 : _T_1035; // @[LZD.scala 49:35]
  assign _T_1038 = {_T_1031,_T_1033,_T_1036}; // @[Cat.scala 29:58]
  assign _T_1039 = _T_1013[2]; // @[Shift.scala 12:21]
  assign _T_1040 = _T_1038[2]; // @[Shift.scala 12:21]
  assign _T_1041 = _T_1039 | _T_1040; // @[LZD.scala 49:16]
  assign _T_1042 = ~ _T_1040; // @[LZD.scala 49:27]
  assign _T_1043 = _T_1039 | _T_1042; // @[LZD.scala 49:25]
  assign _T_1044 = _T_1013[1:0]; // @[LZD.scala 49:47]
  assign _T_1045 = _T_1038[1:0]; // @[LZD.scala 49:59]
  assign _T_1046 = _T_1039 ? _T_1044 : _T_1045; // @[LZD.scala 49:35]
  assign _T_1048 = {_T_1041,_T_1043,_T_1046}; // @[Cat.scala 29:58]
  assign _T_1049 = _T_987[6:0]; // @[LZD.scala 44:32]
  assign _T_1050 = _T_1049[6:3]; // @[LZD.scala 43:32]
  assign _T_1051 = _T_1050[3:2]; // @[LZD.scala 43:32]
  assign _T_1052 = _T_1051 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1053 = _T_1051[1]; // @[LZD.scala 39:21]
  assign _T_1054 = _T_1051[0]; // @[LZD.scala 39:30]
  assign _T_1055 = ~ _T_1054; // @[LZD.scala 39:27]
  assign _T_1056 = _T_1053 | _T_1055; // @[LZD.scala 39:25]
  assign _T_1057 = {_T_1052,_T_1056}; // @[Cat.scala 29:58]
  assign _T_1058 = _T_1050[1:0]; // @[LZD.scala 44:32]
  assign _T_1059 = _T_1058 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1060 = _T_1058[1]; // @[LZD.scala 39:21]
  assign _T_1061 = _T_1058[0]; // @[LZD.scala 39:30]
  assign _T_1062 = ~ _T_1061; // @[LZD.scala 39:27]
  assign _T_1063 = _T_1060 | _T_1062; // @[LZD.scala 39:25]
  assign _T_1064 = {_T_1059,_T_1063}; // @[Cat.scala 29:58]
  assign _T_1065 = _T_1057[1]; // @[Shift.scala 12:21]
  assign _T_1066 = _T_1064[1]; // @[Shift.scala 12:21]
  assign _T_1067 = _T_1065 | _T_1066; // @[LZD.scala 49:16]
  assign _T_1068 = ~ _T_1066; // @[LZD.scala 49:27]
  assign _T_1069 = _T_1065 | _T_1068; // @[LZD.scala 49:25]
  assign _T_1070 = _T_1057[0:0]; // @[LZD.scala 49:47]
  assign _T_1071 = _T_1064[0:0]; // @[LZD.scala 49:59]
  assign _T_1072 = _T_1065 ? _T_1070 : _T_1071; // @[LZD.scala 49:35]
  assign _T_1074 = {_T_1067,_T_1069,_T_1072}; // @[Cat.scala 29:58]
  assign _T_1075 = _T_1049[2:0]; // @[LZD.scala 44:32]
  assign _T_1076 = _T_1075[2:1]; // @[LZD.scala 43:32]
  assign _T_1077 = _T_1076 != 2'h0; // @[LZD.scala 39:14]
  assign _T_1078 = _T_1076[1]; // @[LZD.scala 39:21]
  assign _T_1079 = _T_1076[0]; // @[LZD.scala 39:30]
  assign _T_1080 = ~ _T_1079; // @[LZD.scala 39:27]
  assign _T_1081 = _T_1078 | _T_1080; // @[LZD.scala 39:25]
  assign _T_1082 = {_T_1077,_T_1081}; // @[Cat.scala 29:58]
  assign _T_1083 = _T_1075[0:0]; // @[LZD.scala 44:32]
  assign _T_1085 = _T_1082[1]; // @[Shift.scala 12:21]
  assign _T_1087 = _T_1082[0:0]; // @[LZD.scala 55:32]
  assign _T_1088 = _T_1085 ? _T_1087 : _T_1083; // @[LZD.scala 55:20]
  assign _T_1089 = {_T_1085,_T_1088}; // @[Cat.scala 29:58]
  assign _T_1090 = _T_1074[2]; // @[Shift.scala 12:21]
  assign _T_1092 = _T_1074[1:0]; // @[LZD.scala 55:32]
  assign _T_1093 = _T_1090 ? _T_1092 : _T_1089; // @[LZD.scala 55:20]
  assign _T_1094 = {_T_1090,_T_1093}; // @[Cat.scala 29:58]
  assign _T_1095 = _T_1048[3]; // @[Shift.scala 12:21]
  assign _T_1097 = _T_1048[2:0]; // @[LZD.scala 55:32]
  assign _T_1098 = _T_1095 ? _T_1097 : _T_1094; // @[LZD.scala 55:20]
  assign _T_1099 = {_T_1095,_T_1098}; // @[Cat.scala 29:58]
  assign _T_1100 = _T_986[4]; // @[Shift.scala 12:21]
  assign _T_1102 = _T_986[3:0]; // @[LZD.scala 55:32]
  assign _T_1103 = _T_1100 ? _T_1102 : _T_1099; // @[LZD.scala 55:20]
  assign _T_1104 = {_T_1100,_T_1103}; // @[Cat.scala 29:58]
  assign _T_1105 = _T_852[5]; // @[Shift.scala 12:21]
  assign _T_1107 = _T_852[4:0]; // @[LZD.scala 55:32]
  assign _T_1108 = _T_1105 ? _T_1107 : _T_1104; // @[LZD.scala 55:20]
  assign _T_1109 = {_T_1105,_T_1108}; // @[Cat.scala 29:58]
  assign _T_1110 = _T_574[6]; // @[Shift.scala 12:21]
  assign _T_1112 = _T_574[5:0]; // @[LZD.scala 55:32]
  assign _T_1113 = _T_1110 ? _T_1112 : _T_1109; // @[LZD.scala 55:20]
  assign scaleBias = {1'h1,_T_1110,_T_1113}; // @[Cat.scala 29:58]
  assign _T_1114 = $signed(scaleBias); // @[QuireToPosit.scala 61:53]
  assign _GEN_2 = {{1{_T_1114[7]}},_T_1114}; // @[QuireToPosit.scala 61:41]
  assign _T_1116 = $signed(9'sh4f) + $signed(_GEN_2); // @[QuireToPosit.scala 61:41]
  assign realScale = $signed(_T_1116); // @[QuireToPosit.scala 61:41]
  assign underflow = $signed(realScale) < $signed(-9'sh18); // @[QuireToPosit.scala 62:41]
  assign overflow = $signed(realScale) > $signed(9'sh18); // @[QuireToPosit.scala 63:35]
  assign _T_1117 = underflow ? $signed(-9'sh18) : $signed(realScale); // @[Mux.scala 87:16]
  assign _T_1118 = overflow ? $signed(9'sh18) : $signed(_T_1117); // @[Mux.scala 87:16]
  assign _T_1119 = realScale[8:8]; // @[Abs.scala 10:21]
  assign _T_1121 = _T_1119 ? 9'h1ff : 9'h0; // @[Bitwise.scala 71:12]
  assign _T_1122 = $unsigned(realScale); // @[Abs.scala 10:31]
  assign _T_1123 = _T_1121 ^ _T_1122; // @[Abs.scala 10:26]
  assign _GEN_3 = {{8'd0}, _T_1119}; // @[Abs.scala 10:39]
  assign absRealScale = _T_1123 + _GEN_3; // @[Abs.scala 10:39]
  assign _T_1126 = absRealScale < 9'h80; // @[Shift.scala 16:24]
  assign _T_1127 = absRealScale[6:0]; // @[Shift.scala 17:37]
  assign _T_1128 = _T_1127[6]; // @[Shift.scala 12:21]
  assign _T_1129 = io_quireIn[63:0]; // @[Shift.scala 64:52]
  assign _T_1131 = {_T_1129,64'h0}; // @[Cat.scala 29:58]
  assign _T_1132 = _T_1128 ? _T_1131 : io_quireIn; // @[Shift.scala 64:27]
  assign _T_1133 = _T_1127[5:0]; // @[Shift.scala 66:70]
  assign _T_1134 = _T_1133[5]; // @[Shift.scala 12:21]
  assign _T_1135 = _T_1132[95:0]; // @[Shift.scala 64:52]
  assign _T_1137 = {_T_1135,32'h0}; // @[Cat.scala 29:58]
  assign _T_1138 = _T_1134 ? _T_1137 : _T_1132; // @[Shift.scala 64:27]
  assign _T_1139 = _T_1133[4:0]; // @[Shift.scala 66:70]
  assign _T_1140 = _T_1139[4]; // @[Shift.scala 12:21]
  assign _T_1141 = _T_1138[111:0]; // @[Shift.scala 64:52]
  assign _T_1143 = {_T_1141,16'h0}; // @[Cat.scala 29:58]
  assign _T_1144 = _T_1140 ? _T_1143 : _T_1138; // @[Shift.scala 64:27]
  assign _T_1145 = _T_1139[3:0]; // @[Shift.scala 66:70]
  assign _T_1146 = _T_1145[3]; // @[Shift.scala 12:21]
  assign _T_1147 = _T_1144[119:0]; // @[Shift.scala 64:52]
  assign _T_1149 = {_T_1147,8'h0}; // @[Cat.scala 29:58]
  assign _T_1150 = _T_1146 ? _T_1149 : _T_1144; // @[Shift.scala 64:27]
  assign _T_1151 = _T_1145[2:0]; // @[Shift.scala 66:70]
  assign _T_1152 = _T_1151[2]; // @[Shift.scala 12:21]
  assign _T_1153 = _T_1150[123:0]; // @[Shift.scala 64:52]
  assign _T_1155 = {_T_1153,4'h0}; // @[Cat.scala 29:58]
  assign _T_1156 = _T_1152 ? _T_1155 : _T_1150; // @[Shift.scala 64:27]
  assign _T_1157 = _T_1151[1:0]; // @[Shift.scala 66:70]
  assign _T_1158 = _T_1157[1]; // @[Shift.scala 12:21]
  assign _T_1159 = _T_1156[125:0]; // @[Shift.scala 64:52]
  assign _T_1161 = {_T_1159,2'h0}; // @[Cat.scala 29:58]
  assign _T_1162 = _T_1158 ? _T_1161 : _T_1156; // @[Shift.scala 64:27]
  assign _T_1163 = _T_1157[0:0]; // @[Shift.scala 66:70]
  assign _T_1165 = _T_1162[126:0]; // @[Shift.scala 64:52]
  assign _T_1166 = {_T_1165,1'h0}; // @[Cat.scala 29:58]
  assign _T_1167 = _T_1163 ? _T_1166 : _T_1162; // @[Shift.scala 64:27]
  assign quireLeftShift = _T_1126 ? _T_1167 : 128'h0; // @[Shift.scala 16:10]
  assign _T_1172 = io_quireIn[127:64]; // @[Shift.scala 77:66]
  assign _T_1173 = {64'h0,_T_1172}; // @[Cat.scala 29:58]
  assign _T_1174 = _T_1128 ? _T_1173 : io_quireIn; // @[Shift.scala 77:22]
  assign _T_1178 = _T_1174[127:32]; // @[Shift.scala 77:66]
  assign _T_1179 = {32'h0,_T_1178}; // @[Cat.scala 29:58]
  assign _T_1180 = _T_1134 ? _T_1179 : _T_1174; // @[Shift.scala 77:22]
  assign _T_1184 = _T_1180[127:16]; // @[Shift.scala 77:66]
  assign _T_1185 = {16'h0,_T_1184}; // @[Cat.scala 29:58]
  assign _T_1186 = _T_1140 ? _T_1185 : _T_1180; // @[Shift.scala 77:22]
  assign _T_1190 = _T_1186[127:8]; // @[Shift.scala 77:66]
  assign _T_1191 = {8'h0,_T_1190}; // @[Cat.scala 29:58]
  assign _T_1192 = _T_1146 ? _T_1191 : _T_1186; // @[Shift.scala 77:22]
  assign _T_1196 = _T_1192[127:4]; // @[Shift.scala 77:66]
  assign _T_1197 = {4'h0,_T_1196}; // @[Cat.scala 29:58]
  assign _T_1198 = _T_1152 ? _T_1197 : _T_1192; // @[Shift.scala 77:22]
  assign _T_1202 = _T_1198[127:2]; // @[Shift.scala 77:66]
  assign _T_1203 = {2'h0,_T_1202}; // @[Cat.scala 29:58]
  assign _T_1204 = _T_1158 ? _T_1203 : _T_1198; // @[Shift.scala 77:22]
  assign _T_1207 = _T_1204[127:1]; // @[Shift.scala 77:66]
  assign _T_1208 = {1'h0,_T_1207}; // @[Cat.scala 29:58]
  assign _T_1209 = _T_1163 ? _T_1208 : _T_1204; // @[Shift.scala 77:22]
  assign quireRightShift = _T_1126 ? _T_1209 : 128'h0; // @[Shift.scala 27:10]
  assign _T_1211 = quireLeftShift[47:43]; // @[QuireToPosit.scala 89:49]
  assign _T_1212 = quireLeftShift[42:0]; // @[QuireToPosit.scala 90:127]
  assign _T_1213 = _T_1212 != 43'h0; // @[QuireToPosit.scala 90:154]
  assign realFGRSTmp1 = {_T_1211,_T_1213}; // @[Cat.scala 29:58]
  assign _T_1214 = quireRightShift[47:43]; // @[QuireToPosit.scala 91:50]
  assign _T_1215 = quireRightShift[42:0]; // @[QuireToPosit.scala 92:128]
  assign _T_1216 = _T_1215 != 43'h0; // @[QuireToPosit.scala 92:155]
  assign realFGRSTmp2 = {_T_1214,_T_1216}; // @[Cat.scala 29:58]
  assign realFGRS = _T_1119 ? realFGRSTmp1 : realFGRSTmp2; // @[QuireToPosit.scala 93:34]
  assign outRawFloat_fraction = realFGRS[5:3]; // @[QuireToPosit.scala 95:46]
  assign outRawFloat_grs = realFGRS[2:0]; // @[QuireToPosit.scala 96:46]
  assign _GEN_4 = _T_1118[5:0]; // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign outRawFloat_scale = $signed(_GEN_4); // @[QuireToPosit.scala 44:31 QuireToPosit.scala 65:27]
  assign _T_1221 = outRawFloat_scale[1:0]; // @[convert.scala 46:61]
  assign _T_1222 = ~ _T_1221; // @[convert.scala 46:52]
  assign _T_1224 = _T_2 ? _T_1222 : _T_1221; // @[convert.scala 46:42]
  assign _T_1225 = outRawFloat_scale[5:2]; // @[convert.scala 48:34]
  assign _T_1226 = _T_1225[3:3]; // @[convert.scala 49:36]
  assign _T_1228 = ~ _T_1225; // @[convert.scala 50:36]
  assign _T_1229 = $signed(_T_1228); // @[convert.scala 50:36]
  assign _T_1230 = _T_1226 ? $signed(_T_1229) : $signed(_T_1225); // @[convert.scala 50:28]
  assign _T_1231 = _T_1226 ^ _T_2; // @[convert.scala 51:31]
  assign _T_1232 = ~ _T_1231; // @[convert.scala 52:43]
  assign _T_1236 = {_T_1232,_T_1231,_T_1224,outRawFloat_fraction,outRawFloat_grs}; // @[Cat.scala 29:58]
  assign _T_1237 = $unsigned(_T_1230); // @[Shift.scala 39:17]
  assign _T_1238 = _T_1237 < 4'ha; // @[Shift.scala 39:24]
  assign _T_1240 = _T_1236[9:8]; // @[Shift.scala 90:30]
  assign _T_1241 = _T_1236[7:0]; // @[Shift.scala 90:48]
  assign _T_1242 = _T_1241 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{1'd0}, _T_1242}; // @[Shift.scala 90:39]
  assign _T_1243 = _T_1240 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_1244 = _T_1237[3]; // @[Shift.scala 12:21]
  assign _T_1245 = _T_1236[9]; // @[Shift.scala 12:21]
  assign _T_1247 = _T_1245 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_1248 = {_T_1247,_T_1243}; // @[Cat.scala 29:58]
  assign _T_1249 = _T_1244 ? _T_1248 : _T_1236; // @[Shift.scala 91:22]
  assign _T_1250 = _T_1237[2:0]; // @[Shift.scala 92:77]
  assign _T_1251 = _T_1249[9:4]; // @[Shift.scala 90:30]
  assign _T_1252 = _T_1249[3:0]; // @[Shift.scala 90:48]
  assign _T_1253 = _T_1252 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_6 = {{5'd0}, _T_1253}; // @[Shift.scala 90:39]
  assign _T_1254 = _T_1251 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_1255 = _T_1250[2]; // @[Shift.scala 12:21]
  assign _T_1256 = _T_1249[9]; // @[Shift.scala 12:21]
  assign _T_1258 = _T_1256 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_1259 = {_T_1258,_T_1254}; // @[Cat.scala 29:58]
  assign _T_1260 = _T_1255 ? _T_1259 : _T_1249; // @[Shift.scala 91:22]
  assign _T_1261 = _T_1250[1:0]; // @[Shift.scala 92:77]
  assign _T_1262 = _T_1260[9:2]; // @[Shift.scala 90:30]
  assign _T_1263 = _T_1260[1:0]; // @[Shift.scala 90:48]
  assign _T_1264 = _T_1263 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_7 = {{7'd0}, _T_1264}; // @[Shift.scala 90:39]
  assign _T_1265 = _T_1262 | _GEN_7; // @[Shift.scala 90:39]
  assign _T_1266 = _T_1261[1]; // @[Shift.scala 12:21]
  assign _T_1267 = _T_1260[9]; // @[Shift.scala 12:21]
  assign _T_1269 = _T_1267 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_1270 = {_T_1269,_T_1265}; // @[Cat.scala 29:58]
  assign _T_1271 = _T_1266 ? _T_1270 : _T_1260; // @[Shift.scala 91:22]
  assign _T_1272 = _T_1261[0:0]; // @[Shift.scala 92:77]
  assign _T_1273 = _T_1271[9:1]; // @[Shift.scala 90:30]
  assign _T_1274 = _T_1271[0:0]; // @[Shift.scala 90:48]
  assign _GEN_8 = {{8'd0}, _T_1274}; // @[Shift.scala 90:39]
  assign _T_1276 = _T_1273 | _GEN_8; // @[Shift.scala 90:39]
  assign _T_1278 = _T_1271[9]; // @[Shift.scala 12:21]
  assign _T_1279 = {_T_1278,_T_1276}; // @[Cat.scala 29:58]
  assign _T_1280 = _T_1272 ? _T_1279 : _T_1271; // @[Shift.scala 91:22]
  assign _T_1283 = _T_1245 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign _T_1284 = _T_1238 ? _T_1280 : _T_1283; // @[Shift.scala 39:10]
  assign _T_1285 = _T_1284[3]; // @[convert.scala 55:31]
  assign _T_1286 = _T_1284[2]; // @[convert.scala 56:31]
  assign _T_1287 = _T_1284[1]; // @[convert.scala 57:31]
  assign _T_1288 = _T_1284[0]; // @[convert.scala 58:31]
  assign _T_1289 = _T_1284[9:3]; // @[convert.scala 59:69]
  assign _T_1290 = _T_1289 != 7'h0; // @[convert.scala 59:81]
  assign _T_1291 = ~ _T_1290; // @[convert.scala 59:50]
  assign _T_1293 = _T_1289 == 7'h7f; // @[convert.scala 60:81]
  assign _T_1294 = _T_1285 | _T_1287; // @[convert.scala 61:44]
  assign _T_1295 = _T_1294 | _T_1288; // @[convert.scala 61:52]
  assign _T_1296 = _T_1286 & _T_1295; // @[convert.scala 61:36]
  assign _T_1297 = ~ _T_1293; // @[convert.scala 62:63]
  assign _T_1298 = _T_1297 & _T_1296; // @[convert.scala 62:103]
  assign _T_1299 = _T_1291 | _T_1298; // @[convert.scala 62:60]
  assign _GEN_9 = {{6'd0}, _T_1299}; // @[convert.scala 63:56]
  assign _T_1302 = _T_1289 + _GEN_9; // @[convert.scala 63:56]
  assign _T_1303 = {_T_2,_T_1302}; // @[Cat.scala 29:58]
  assign io_positOut = _T_1311; // @[QuireToPosit.scala 101:15]
  assign io_outValid = _T_1307; // @[QuireToPosit.scala 100:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1307 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1311 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      _T_1307 <= 1'h0;
    end else begin
      _T_1307 <= io_inValid;
    end
    if (io_inValid) begin
      if (outRawFloat_isNaR) begin
        _T_1311 <= 8'h80;
      end else begin
        if (outRawFloat_isZero) begin
          _T_1311 <= 8'h0;
        end else begin
          _T_1311 <= _T_1303;
        end
      end
    end
  end
endmodule
