module PositMultiplier16_4(
  input         clock,
  input         reset,
  input  [15:0] io_A,
  input  [15:0] io_B,
  output [15:0] io_M
);
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [13:0] _T_4; // @[convert.scala 19:24]
  wire [13:0] _T_5; // @[convert.scala 19:43]
  wire [13:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [5:0] _T_68; // @[LZD.scala 44:32]
  wire [3:0] _T_69; // @[LZD.scala 43:32]
  wire [1:0] _T_70; // @[LZD.scala 43:32]
  wire  _T_71; // @[LZD.scala 39:14]
  wire  _T_72; // @[LZD.scala 39:21]
  wire  _T_73; // @[LZD.scala 39:30]
  wire  _T_74; // @[LZD.scala 39:27]
  wire  _T_75; // @[LZD.scala 39:25]
  wire [1:0] _T_76; // @[Cat.scala 29:58]
  wire [1:0] _T_77; // @[LZD.scala 44:32]
  wire  _T_78; // @[LZD.scala 39:14]
  wire  _T_79; // @[LZD.scala 39:21]
  wire  _T_80; // @[LZD.scala 39:30]
  wire  _T_81; // @[LZD.scala 39:27]
  wire  _T_82; // @[LZD.scala 39:25]
  wire [1:0] _T_83; // @[Cat.scala 29:58]
  wire  _T_84; // @[Shift.scala 12:21]
  wire  _T_85; // @[Shift.scala 12:21]
  wire  _T_86; // @[LZD.scala 49:16]
  wire  _T_87; // @[LZD.scala 49:27]
  wire  _T_88; // @[LZD.scala 49:25]
  wire  _T_89; // @[LZD.scala 49:47]
  wire  _T_90; // @[LZD.scala 49:59]
  wire  _T_91; // @[LZD.scala 49:35]
  wire [2:0] _T_93; // @[Cat.scala 29:58]
  wire [1:0] _T_94; // @[LZD.scala 44:32]
  wire  _T_95; // @[LZD.scala 39:14]
  wire  _T_96; // @[LZD.scala 39:21]
  wire  _T_97; // @[LZD.scala 39:30]
  wire  _T_98; // @[LZD.scala 39:27]
  wire  _T_99; // @[LZD.scala 39:25]
  wire [1:0] _T_100; // @[Cat.scala 29:58]
  wire  _T_101; // @[Shift.scala 12:21]
  wire [1:0] _T_103; // @[LZD.scala 55:32]
  wire [1:0] _T_104; // @[LZD.scala 55:20]
  wire [2:0] _T_105; // @[Cat.scala 29:58]
  wire  _T_106; // @[Shift.scala 12:21]
  wire [2:0] _T_108; // @[LZD.scala 55:32]
  wire [2:0] _T_109; // @[LZD.scala 55:20]
  wire [3:0] _T_110; // @[Cat.scala 29:58]
  wire [3:0] _T_111; // @[convert.scala 21:22]
  wire [12:0] _T_112; // @[convert.scala 22:36]
  wire  _T_113; // @[Shift.scala 16:24]
  wire  _T_115; // @[Shift.scala 12:21]
  wire [4:0] _T_116; // @[Shift.scala 64:52]
  wire [12:0] _T_118; // @[Cat.scala 29:58]
  wire [12:0] _T_119; // @[Shift.scala 64:27]
  wire [2:0] _T_120; // @[Shift.scala 66:70]
  wire  _T_121; // @[Shift.scala 12:21]
  wire [8:0] _T_122; // @[Shift.scala 64:52]
  wire [12:0] _T_124; // @[Cat.scala 29:58]
  wire [12:0] _T_125; // @[Shift.scala 64:27]
  wire [1:0] _T_126; // @[Shift.scala 66:70]
  wire  _T_127; // @[Shift.scala 12:21]
  wire [10:0] _T_128; // @[Shift.scala 64:52]
  wire [12:0] _T_130; // @[Cat.scala 29:58]
  wire [12:0] _T_131; // @[Shift.scala 64:27]
  wire  _T_132; // @[Shift.scala 66:70]
  wire [11:0] _T_134; // @[Shift.scala 64:52]
  wire [12:0] _T_135; // @[Cat.scala 29:58]
  wire [12:0] _T_136; // @[Shift.scala 64:27]
  wire [12:0] _T_137; // @[Shift.scala 16:10]
  wire [3:0] _T_138; // @[convert.scala 23:34]
  wire [8:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_140; // @[convert.scala 25:26]
  wire [3:0] _T_142; // @[convert.scala 25:42]
  wire [3:0] _T_145; // @[convert.scala 26:67]
  wire [3:0] _T_146; // @[convert.scala 26:51]
  wire [8:0] _T_147; // @[Cat.scala 29:58]
  wire [14:0] _T_149; // @[convert.scala 29:56]
  wire  _T_150; // @[convert.scala 29:60]
  wire  _T_151; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_154; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [8:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_163; // @[convert.scala 18:24]
  wire  _T_164; // @[convert.scala 18:40]
  wire  _T_165; // @[convert.scala 18:36]
  wire [13:0] _T_166; // @[convert.scala 19:24]
  wire [13:0] _T_167; // @[convert.scala 19:43]
  wire [13:0] _T_168; // @[convert.scala 19:39]
  wire [7:0] _T_169; // @[LZD.scala 43:32]
  wire [3:0] _T_170; // @[LZD.scala 43:32]
  wire [1:0] _T_171; // @[LZD.scala 43:32]
  wire  _T_172; // @[LZD.scala 39:14]
  wire  _T_173; // @[LZD.scala 39:21]
  wire  _T_174; // @[LZD.scala 39:30]
  wire  _T_175; // @[LZD.scala 39:27]
  wire  _T_176; // @[LZD.scala 39:25]
  wire [1:0] _T_177; // @[Cat.scala 29:58]
  wire [1:0] _T_178; // @[LZD.scala 44:32]
  wire  _T_179; // @[LZD.scala 39:14]
  wire  _T_180; // @[LZD.scala 39:21]
  wire  _T_181; // @[LZD.scala 39:30]
  wire  _T_182; // @[LZD.scala 39:27]
  wire  _T_183; // @[LZD.scala 39:25]
  wire [1:0] _T_184; // @[Cat.scala 29:58]
  wire  _T_185; // @[Shift.scala 12:21]
  wire  _T_186; // @[Shift.scala 12:21]
  wire  _T_187; // @[LZD.scala 49:16]
  wire  _T_188; // @[LZD.scala 49:27]
  wire  _T_189; // @[LZD.scala 49:25]
  wire  _T_190; // @[LZD.scala 49:47]
  wire  _T_191; // @[LZD.scala 49:59]
  wire  _T_192; // @[LZD.scala 49:35]
  wire [2:0] _T_194; // @[Cat.scala 29:58]
  wire [3:0] _T_195; // @[LZD.scala 44:32]
  wire [1:0] _T_196; // @[LZD.scala 43:32]
  wire  _T_197; // @[LZD.scala 39:14]
  wire  _T_198; // @[LZD.scala 39:21]
  wire  _T_199; // @[LZD.scala 39:30]
  wire  _T_200; // @[LZD.scala 39:27]
  wire  _T_201; // @[LZD.scala 39:25]
  wire [1:0] _T_202; // @[Cat.scala 29:58]
  wire [1:0] _T_203; // @[LZD.scala 44:32]
  wire  _T_204; // @[LZD.scala 39:14]
  wire  _T_205; // @[LZD.scala 39:21]
  wire  _T_206; // @[LZD.scala 39:30]
  wire  _T_207; // @[LZD.scala 39:27]
  wire  _T_208; // @[LZD.scala 39:25]
  wire [1:0] _T_209; // @[Cat.scala 29:58]
  wire  _T_210; // @[Shift.scala 12:21]
  wire  _T_211; // @[Shift.scala 12:21]
  wire  _T_212; // @[LZD.scala 49:16]
  wire  _T_213; // @[LZD.scala 49:27]
  wire  _T_214; // @[LZD.scala 49:25]
  wire  _T_215; // @[LZD.scala 49:47]
  wire  _T_216; // @[LZD.scala 49:59]
  wire  _T_217; // @[LZD.scala 49:35]
  wire [2:0] _T_219; // @[Cat.scala 29:58]
  wire  _T_220; // @[Shift.scala 12:21]
  wire  _T_221; // @[Shift.scala 12:21]
  wire  _T_222; // @[LZD.scala 49:16]
  wire  _T_223; // @[LZD.scala 49:27]
  wire  _T_224; // @[LZD.scala 49:25]
  wire [1:0] _T_225; // @[LZD.scala 49:47]
  wire [1:0] _T_226; // @[LZD.scala 49:59]
  wire [1:0] _T_227; // @[LZD.scala 49:35]
  wire [3:0] _T_229; // @[Cat.scala 29:58]
  wire [5:0] _T_230; // @[LZD.scala 44:32]
  wire [3:0] _T_231; // @[LZD.scala 43:32]
  wire [1:0] _T_232; // @[LZD.scala 43:32]
  wire  _T_233; // @[LZD.scala 39:14]
  wire  _T_234; // @[LZD.scala 39:21]
  wire  _T_235; // @[LZD.scala 39:30]
  wire  _T_236; // @[LZD.scala 39:27]
  wire  _T_237; // @[LZD.scala 39:25]
  wire [1:0] _T_238; // @[Cat.scala 29:58]
  wire [1:0] _T_239; // @[LZD.scala 44:32]
  wire  _T_240; // @[LZD.scala 39:14]
  wire  _T_241; // @[LZD.scala 39:21]
  wire  _T_242; // @[LZD.scala 39:30]
  wire  _T_243; // @[LZD.scala 39:27]
  wire  _T_244; // @[LZD.scala 39:25]
  wire [1:0] _T_245; // @[Cat.scala 29:58]
  wire  _T_246; // @[Shift.scala 12:21]
  wire  _T_247; // @[Shift.scala 12:21]
  wire  _T_248; // @[LZD.scala 49:16]
  wire  _T_249; // @[LZD.scala 49:27]
  wire  _T_250; // @[LZD.scala 49:25]
  wire  _T_251; // @[LZD.scala 49:47]
  wire  _T_252; // @[LZD.scala 49:59]
  wire  _T_253; // @[LZD.scala 49:35]
  wire [2:0] _T_255; // @[Cat.scala 29:58]
  wire [1:0] _T_256; // @[LZD.scala 44:32]
  wire  _T_257; // @[LZD.scala 39:14]
  wire  _T_258; // @[LZD.scala 39:21]
  wire  _T_259; // @[LZD.scala 39:30]
  wire  _T_260; // @[LZD.scala 39:27]
  wire  _T_261; // @[LZD.scala 39:25]
  wire [1:0] _T_262; // @[Cat.scala 29:58]
  wire  _T_263; // @[Shift.scala 12:21]
  wire [1:0] _T_265; // @[LZD.scala 55:32]
  wire [1:0] _T_266; // @[LZD.scala 55:20]
  wire [2:0] _T_267; // @[Cat.scala 29:58]
  wire  _T_268; // @[Shift.scala 12:21]
  wire [2:0] _T_270; // @[LZD.scala 55:32]
  wire [2:0] _T_271; // @[LZD.scala 55:20]
  wire [3:0] _T_272; // @[Cat.scala 29:58]
  wire [3:0] _T_273; // @[convert.scala 21:22]
  wire [12:0] _T_274; // @[convert.scala 22:36]
  wire  _T_275; // @[Shift.scala 16:24]
  wire  _T_277; // @[Shift.scala 12:21]
  wire [4:0] _T_278; // @[Shift.scala 64:52]
  wire [12:0] _T_280; // @[Cat.scala 29:58]
  wire [12:0] _T_281; // @[Shift.scala 64:27]
  wire [2:0] _T_282; // @[Shift.scala 66:70]
  wire  _T_283; // @[Shift.scala 12:21]
  wire [8:0] _T_284; // @[Shift.scala 64:52]
  wire [12:0] _T_286; // @[Cat.scala 29:58]
  wire [12:0] _T_287; // @[Shift.scala 64:27]
  wire [1:0] _T_288; // @[Shift.scala 66:70]
  wire  _T_289; // @[Shift.scala 12:21]
  wire [10:0] _T_290; // @[Shift.scala 64:52]
  wire [12:0] _T_292; // @[Cat.scala 29:58]
  wire [12:0] _T_293; // @[Shift.scala 64:27]
  wire  _T_294; // @[Shift.scala 66:70]
  wire [11:0] _T_296; // @[Shift.scala 64:52]
  wire [12:0] _T_297; // @[Cat.scala 29:58]
  wire [12:0] _T_298; // @[Shift.scala 64:27]
  wire [12:0] _T_299; // @[Shift.scala 16:10]
  wire [3:0] _T_300; // @[convert.scala 23:34]
  wire [8:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_302; // @[convert.scala 25:26]
  wire [3:0] _T_304; // @[convert.scala 25:42]
  wire [3:0] _T_307; // @[convert.scala 26:67]
  wire [3:0] _T_308; // @[convert.scala 26:51]
  wire [8:0] _T_309; // @[Cat.scala 29:58]
  wire [14:0] _T_311; // @[convert.scala 29:56]
  wire  _T_312; // @[convert.scala 29:60]
  wire  _T_313; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_316; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [8:0] decB_scale; // @[convert.scala 32:24]
  wire  _T_324; // @[PositMultiplier.scala 43:34]
  wire [10:0] _T_326; // @[Cat.scala 29:58]
  wire [10:0] sigA; // @[PositMultiplier.scala 43:61]
  wire  _T_327; // @[PositMultiplier.scala 44:34]
  wire [10:0] _T_329; // @[Cat.scala 29:58]
  wire [10:0] sigB; // @[PositMultiplier.scala 44:61]
  wire [21:0] _T_330; // @[PositMultiplier.scala 45:25]
  wire [21:0] sigP; // @[PositMultiplier.scala 45:33]
  wire [1:0] head2; // @[PositMultiplier.scala 46:28]
  wire  _T_331; // @[PositMultiplier.scala 47:31]
  wire  _T_332; // @[PositMultiplier.scala 47:25]
  wire  _T_333; // @[PositMultiplier.scala 47:42]
  wire  addTwo; // @[PositMultiplier.scala 47:35]
  wire  _T_334; // @[PositMultiplier.scala 49:23]
  wire  _T_335; // @[PositMultiplier.scala 49:49]
  wire  addOne; // @[PositMultiplier.scala 49:43]
  wire [1:0] _T_336; // @[Cat.scala 29:58]
  wire [2:0] expBias; // @[PositMultiplier.scala 50:39]
  wire [18:0] _T_337; // @[PositMultiplier.scala 53:81]
  wire [17:0] _T_338; // @[PositMultiplier.scala 54:81]
  wire [18:0] _T_339; // @[PositMultiplier.scala 54:104]
  wire [18:0] frac; // @[PositMultiplier.scala 51:22]
  wire [9:0] _T_340; // @[PositMultiplier.scala 56:30]
  wire [9:0] _GEN_0; // @[PositMultiplier.scala 56:44]
  wire [9:0] _T_342; // @[PositMultiplier.scala 56:44]
  wire [9:0] mulScale; // @[PositMultiplier.scala 56:44]
  wire  underflow; // @[PositMultiplier.scala 57:28]
  wire  overflow; // @[PositMultiplier.scala 58:28]
  wire  decM_sign; // @[PositMultiplier.scala 62:29]
  wire [9:0] _T_345; // @[Mux.scala 87:16]
  wire [9:0] _T_346; // @[Mux.scala 87:16]
  wire [8:0] decM_fraction; // @[PositMultiplier.scala 70:29]
  wire  decM_isNaR; // @[PositMultiplier.scala 71:31]
  wire  decM_isZero; // @[PositMultiplier.scala 72:32]
  wire [9:0] grsTmp; // @[PositMultiplier.scala 75:30]
  wire [1:0] _T_350; // @[PositMultiplier.scala 78:32]
  wire [7:0] _T_351; // @[PositMultiplier.scala 78:48]
  wire  _T_352; // @[PositMultiplier.scala 78:52]
  wire [8:0] _GEN_1; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  wire [8:0] decM_scale; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  wire [3:0] _T_355; // @[convert.scala 46:61]
  wire [3:0] _T_356; // @[convert.scala 46:52]
  wire [3:0] _T_358; // @[convert.scala 46:42]
  wire [4:0] _T_359; // @[convert.scala 48:34]
  wire  _T_360; // @[convert.scala 49:36]
  wire [4:0] _T_362; // @[convert.scala 50:36]
  wire [4:0] _T_363; // @[convert.scala 50:36]
  wire [4:0] _T_364; // @[convert.scala 50:28]
  wire  _T_365; // @[convert.scala 51:31]
  wire  _T_366; // @[convert.scala 52:43]
  wire [17:0] _T_370; // @[Cat.scala 29:58]
  wire [4:0] _T_371; // @[Shift.scala 39:17]
  wire  _T_372; // @[Shift.scala 39:24]
  wire [1:0] _T_374; // @[Shift.scala 90:30]
  wire [15:0] _T_375; // @[Shift.scala 90:48]
  wire  _T_376; // @[Shift.scala 90:57]
  wire [1:0] _GEN_2; // @[Shift.scala 90:39]
  wire [1:0] _T_377; // @[Shift.scala 90:39]
  wire  _T_378; // @[Shift.scala 12:21]
  wire  _T_379; // @[Shift.scala 12:21]
  wire [15:0] _T_381; // @[Bitwise.scala 71:12]
  wire [17:0] _T_382; // @[Cat.scala 29:58]
  wire [17:0] _T_383; // @[Shift.scala 91:22]
  wire [3:0] _T_384; // @[Shift.scala 92:77]
  wire [9:0] _T_385; // @[Shift.scala 90:30]
  wire [7:0] _T_386; // @[Shift.scala 90:48]
  wire  _T_387; // @[Shift.scala 90:57]
  wire [9:0] _GEN_3; // @[Shift.scala 90:39]
  wire [9:0] _T_388; // @[Shift.scala 90:39]
  wire  _T_389; // @[Shift.scala 12:21]
  wire  _T_390; // @[Shift.scala 12:21]
  wire [7:0] _T_392; // @[Bitwise.scala 71:12]
  wire [17:0] _T_393; // @[Cat.scala 29:58]
  wire [17:0] _T_394; // @[Shift.scala 91:22]
  wire [2:0] _T_395; // @[Shift.scala 92:77]
  wire [13:0] _T_396; // @[Shift.scala 90:30]
  wire [3:0] _T_397; // @[Shift.scala 90:48]
  wire  _T_398; // @[Shift.scala 90:57]
  wire [13:0] _GEN_4; // @[Shift.scala 90:39]
  wire [13:0] _T_399; // @[Shift.scala 90:39]
  wire  _T_400; // @[Shift.scala 12:21]
  wire  _T_401; // @[Shift.scala 12:21]
  wire [3:0] _T_403; // @[Bitwise.scala 71:12]
  wire [17:0] _T_404; // @[Cat.scala 29:58]
  wire [17:0] _T_405; // @[Shift.scala 91:22]
  wire [1:0] _T_406; // @[Shift.scala 92:77]
  wire [15:0] _T_407; // @[Shift.scala 90:30]
  wire [1:0] _T_408; // @[Shift.scala 90:48]
  wire  _T_409; // @[Shift.scala 90:57]
  wire [15:0] _GEN_5; // @[Shift.scala 90:39]
  wire [15:0] _T_410; // @[Shift.scala 90:39]
  wire  _T_411; // @[Shift.scala 12:21]
  wire  _T_412; // @[Shift.scala 12:21]
  wire [1:0] _T_414; // @[Bitwise.scala 71:12]
  wire [17:0] _T_415; // @[Cat.scala 29:58]
  wire [17:0] _T_416; // @[Shift.scala 91:22]
  wire  _T_417; // @[Shift.scala 92:77]
  wire [16:0] _T_418; // @[Shift.scala 90:30]
  wire  _T_419; // @[Shift.scala 90:48]
  wire [16:0] _GEN_6; // @[Shift.scala 90:39]
  wire [16:0] _T_421; // @[Shift.scala 90:39]
  wire  _T_423; // @[Shift.scala 12:21]
  wire [17:0] _T_424; // @[Cat.scala 29:58]
  wire [17:0] _T_425; // @[Shift.scala 91:22]
  wire [17:0] _T_428; // @[Bitwise.scala 71:12]
  wire [17:0] _T_429; // @[Shift.scala 39:10]
  wire  _T_430; // @[convert.scala 55:31]
  wire  _T_431; // @[convert.scala 56:31]
  wire  _T_432; // @[convert.scala 57:31]
  wire  _T_433; // @[convert.scala 58:31]
  wire [14:0] _T_434; // @[convert.scala 59:69]
  wire  _T_435; // @[convert.scala 59:81]
  wire  _T_436; // @[convert.scala 59:50]
  wire  _T_438; // @[convert.scala 60:81]
  wire  _T_439; // @[convert.scala 61:44]
  wire  _T_440; // @[convert.scala 61:52]
  wire  _T_441; // @[convert.scala 61:36]
  wire  _T_442; // @[convert.scala 62:63]
  wire  _T_443; // @[convert.scala 62:103]
  wire  _T_444; // @[convert.scala 62:60]
  wire [14:0] _GEN_7; // @[convert.scala 63:56]
  wire [14:0] _T_447; // @[convert.scala 63:56]
  wire [15:0] _T_448; // @[Cat.scala 29:58]
  wire [15:0] _T_450; // @[Mux.scala 87:16]
  assign _T_1 = io_A[15]; // @[convert.scala 18:24]
  assign _T_2 = io_A[14]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[14:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[13:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[13:6]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[5:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68[5:2]; // @[LZD.scala 43:32]
  assign _T_70 = _T_69[3:2]; // @[LZD.scala 43:32]
  assign _T_71 = _T_70 != 2'h0; // @[LZD.scala 39:14]
  assign _T_72 = _T_70[1]; // @[LZD.scala 39:21]
  assign _T_73 = _T_70[0]; // @[LZD.scala 39:30]
  assign _T_74 = ~ _T_73; // @[LZD.scala 39:27]
  assign _T_75 = _T_72 | _T_74; // @[LZD.scala 39:25]
  assign _T_76 = {_T_71,_T_75}; // @[Cat.scala 29:58]
  assign _T_77 = _T_69[1:0]; // @[LZD.scala 44:32]
  assign _T_78 = _T_77 != 2'h0; // @[LZD.scala 39:14]
  assign _T_79 = _T_77[1]; // @[LZD.scala 39:21]
  assign _T_80 = _T_77[0]; // @[LZD.scala 39:30]
  assign _T_81 = ~ _T_80; // @[LZD.scala 39:27]
  assign _T_82 = _T_79 | _T_81; // @[LZD.scala 39:25]
  assign _T_83 = {_T_78,_T_82}; // @[Cat.scala 29:58]
  assign _T_84 = _T_76[1]; // @[Shift.scala 12:21]
  assign _T_85 = _T_83[1]; // @[Shift.scala 12:21]
  assign _T_86 = _T_84 | _T_85; // @[LZD.scala 49:16]
  assign _T_87 = ~ _T_85; // @[LZD.scala 49:27]
  assign _T_88 = _T_84 | _T_87; // @[LZD.scala 49:25]
  assign _T_89 = _T_76[0:0]; // @[LZD.scala 49:47]
  assign _T_90 = _T_83[0:0]; // @[LZD.scala 49:59]
  assign _T_91 = _T_84 ? _T_89 : _T_90; // @[LZD.scala 49:35]
  assign _T_93 = {_T_86,_T_88,_T_91}; // @[Cat.scala 29:58]
  assign _T_94 = _T_68[1:0]; // @[LZD.scala 44:32]
  assign _T_95 = _T_94 != 2'h0; // @[LZD.scala 39:14]
  assign _T_96 = _T_94[1]; // @[LZD.scala 39:21]
  assign _T_97 = _T_94[0]; // @[LZD.scala 39:30]
  assign _T_98 = ~ _T_97; // @[LZD.scala 39:27]
  assign _T_99 = _T_96 | _T_98; // @[LZD.scala 39:25]
  assign _T_100 = {_T_95,_T_99}; // @[Cat.scala 29:58]
  assign _T_101 = _T_93[2]; // @[Shift.scala 12:21]
  assign _T_103 = _T_93[1:0]; // @[LZD.scala 55:32]
  assign _T_104 = _T_101 ? _T_103 : _T_100; // @[LZD.scala 55:20]
  assign _T_105 = {_T_101,_T_104}; // @[Cat.scala 29:58]
  assign _T_106 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_108 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_109 = _T_106 ? _T_108 : _T_105; // @[LZD.scala 55:20]
  assign _T_110 = {_T_106,_T_109}; // @[Cat.scala 29:58]
  assign _T_111 = ~ _T_110; // @[convert.scala 21:22]
  assign _T_112 = io_A[12:0]; // @[convert.scala 22:36]
  assign _T_113 = _T_111 < 4'hd; // @[Shift.scala 16:24]
  assign _T_115 = _T_111[3]; // @[Shift.scala 12:21]
  assign _T_116 = _T_112[4:0]; // @[Shift.scala 64:52]
  assign _T_118 = {_T_116,8'h0}; // @[Cat.scala 29:58]
  assign _T_119 = _T_115 ? _T_118 : _T_112; // @[Shift.scala 64:27]
  assign _T_120 = _T_111[2:0]; // @[Shift.scala 66:70]
  assign _T_121 = _T_120[2]; // @[Shift.scala 12:21]
  assign _T_122 = _T_119[8:0]; // @[Shift.scala 64:52]
  assign _T_124 = {_T_122,4'h0}; // @[Cat.scala 29:58]
  assign _T_125 = _T_121 ? _T_124 : _T_119; // @[Shift.scala 64:27]
  assign _T_126 = _T_120[1:0]; // @[Shift.scala 66:70]
  assign _T_127 = _T_126[1]; // @[Shift.scala 12:21]
  assign _T_128 = _T_125[10:0]; // @[Shift.scala 64:52]
  assign _T_130 = {_T_128,2'h0}; // @[Cat.scala 29:58]
  assign _T_131 = _T_127 ? _T_130 : _T_125; // @[Shift.scala 64:27]
  assign _T_132 = _T_126[0:0]; // @[Shift.scala 66:70]
  assign _T_134 = _T_131[11:0]; // @[Shift.scala 64:52]
  assign _T_135 = {_T_134,1'h0}; // @[Cat.scala 29:58]
  assign _T_136 = _T_132 ? _T_135 : _T_131; // @[Shift.scala 64:27]
  assign _T_137 = _T_113 ? _T_136 : 13'h0; // @[Shift.scala 16:10]
  assign _T_138 = _T_137[12:9]; // @[convert.scala 23:34]
  assign decA_fraction = _T_137[8:0]; // @[convert.scala 24:34]
  assign _T_140 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_142 = _T_3 ? _T_111 : _T_110; // @[convert.scala 25:42]
  assign _T_145 = ~ _T_138; // @[convert.scala 26:67]
  assign _T_146 = _T_1 ? _T_145 : _T_138; // @[convert.scala 26:51]
  assign _T_147 = {_T_140,_T_142,_T_146}; // @[Cat.scala 29:58]
  assign _T_149 = io_A[14:0]; // @[convert.scala 29:56]
  assign _T_150 = _T_149 != 15'h0; // @[convert.scala 29:60]
  assign _T_151 = ~ _T_150; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_151; // @[convert.scala 29:39]
  assign _T_154 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_154 & _T_151; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_147); // @[convert.scala 32:24]
  assign _T_163 = io_B[15]; // @[convert.scala 18:24]
  assign _T_164 = io_B[14]; // @[convert.scala 18:40]
  assign _T_165 = _T_163 ^ _T_164; // @[convert.scala 18:36]
  assign _T_166 = io_B[14:1]; // @[convert.scala 19:24]
  assign _T_167 = io_B[13:0]; // @[convert.scala 19:43]
  assign _T_168 = _T_166 ^ _T_167; // @[convert.scala 19:39]
  assign _T_169 = _T_168[13:6]; // @[LZD.scala 43:32]
  assign _T_170 = _T_169[7:4]; // @[LZD.scala 43:32]
  assign _T_171 = _T_170[3:2]; // @[LZD.scala 43:32]
  assign _T_172 = _T_171 != 2'h0; // @[LZD.scala 39:14]
  assign _T_173 = _T_171[1]; // @[LZD.scala 39:21]
  assign _T_174 = _T_171[0]; // @[LZD.scala 39:30]
  assign _T_175 = ~ _T_174; // @[LZD.scala 39:27]
  assign _T_176 = _T_173 | _T_175; // @[LZD.scala 39:25]
  assign _T_177 = {_T_172,_T_176}; // @[Cat.scala 29:58]
  assign _T_178 = _T_170[1:0]; // @[LZD.scala 44:32]
  assign _T_179 = _T_178 != 2'h0; // @[LZD.scala 39:14]
  assign _T_180 = _T_178[1]; // @[LZD.scala 39:21]
  assign _T_181 = _T_178[0]; // @[LZD.scala 39:30]
  assign _T_182 = ~ _T_181; // @[LZD.scala 39:27]
  assign _T_183 = _T_180 | _T_182; // @[LZD.scala 39:25]
  assign _T_184 = {_T_179,_T_183}; // @[Cat.scala 29:58]
  assign _T_185 = _T_177[1]; // @[Shift.scala 12:21]
  assign _T_186 = _T_184[1]; // @[Shift.scala 12:21]
  assign _T_187 = _T_185 | _T_186; // @[LZD.scala 49:16]
  assign _T_188 = ~ _T_186; // @[LZD.scala 49:27]
  assign _T_189 = _T_185 | _T_188; // @[LZD.scala 49:25]
  assign _T_190 = _T_177[0:0]; // @[LZD.scala 49:47]
  assign _T_191 = _T_184[0:0]; // @[LZD.scala 49:59]
  assign _T_192 = _T_185 ? _T_190 : _T_191; // @[LZD.scala 49:35]
  assign _T_194 = {_T_187,_T_189,_T_192}; // @[Cat.scala 29:58]
  assign _T_195 = _T_169[3:0]; // @[LZD.scala 44:32]
  assign _T_196 = _T_195[3:2]; // @[LZD.scala 43:32]
  assign _T_197 = _T_196 != 2'h0; // @[LZD.scala 39:14]
  assign _T_198 = _T_196[1]; // @[LZD.scala 39:21]
  assign _T_199 = _T_196[0]; // @[LZD.scala 39:30]
  assign _T_200 = ~ _T_199; // @[LZD.scala 39:27]
  assign _T_201 = _T_198 | _T_200; // @[LZD.scala 39:25]
  assign _T_202 = {_T_197,_T_201}; // @[Cat.scala 29:58]
  assign _T_203 = _T_195[1:0]; // @[LZD.scala 44:32]
  assign _T_204 = _T_203 != 2'h0; // @[LZD.scala 39:14]
  assign _T_205 = _T_203[1]; // @[LZD.scala 39:21]
  assign _T_206 = _T_203[0]; // @[LZD.scala 39:30]
  assign _T_207 = ~ _T_206; // @[LZD.scala 39:27]
  assign _T_208 = _T_205 | _T_207; // @[LZD.scala 39:25]
  assign _T_209 = {_T_204,_T_208}; // @[Cat.scala 29:58]
  assign _T_210 = _T_202[1]; // @[Shift.scala 12:21]
  assign _T_211 = _T_209[1]; // @[Shift.scala 12:21]
  assign _T_212 = _T_210 | _T_211; // @[LZD.scala 49:16]
  assign _T_213 = ~ _T_211; // @[LZD.scala 49:27]
  assign _T_214 = _T_210 | _T_213; // @[LZD.scala 49:25]
  assign _T_215 = _T_202[0:0]; // @[LZD.scala 49:47]
  assign _T_216 = _T_209[0:0]; // @[LZD.scala 49:59]
  assign _T_217 = _T_210 ? _T_215 : _T_216; // @[LZD.scala 49:35]
  assign _T_219 = {_T_212,_T_214,_T_217}; // @[Cat.scala 29:58]
  assign _T_220 = _T_194[2]; // @[Shift.scala 12:21]
  assign _T_221 = _T_219[2]; // @[Shift.scala 12:21]
  assign _T_222 = _T_220 | _T_221; // @[LZD.scala 49:16]
  assign _T_223 = ~ _T_221; // @[LZD.scala 49:27]
  assign _T_224 = _T_220 | _T_223; // @[LZD.scala 49:25]
  assign _T_225 = _T_194[1:0]; // @[LZD.scala 49:47]
  assign _T_226 = _T_219[1:0]; // @[LZD.scala 49:59]
  assign _T_227 = _T_220 ? _T_225 : _T_226; // @[LZD.scala 49:35]
  assign _T_229 = {_T_222,_T_224,_T_227}; // @[Cat.scala 29:58]
  assign _T_230 = _T_168[5:0]; // @[LZD.scala 44:32]
  assign _T_231 = _T_230[5:2]; // @[LZD.scala 43:32]
  assign _T_232 = _T_231[3:2]; // @[LZD.scala 43:32]
  assign _T_233 = _T_232 != 2'h0; // @[LZD.scala 39:14]
  assign _T_234 = _T_232[1]; // @[LZD.scala 39:21]
  assign _T_235 = _T_232[0]; // @[LZD.scala 39:30]
  assign _T_236 = ~ _T_235; // @[LZD.scala 39:27]
  assign _T_237 = _T_234 | _T_236; // @[LZD.scala 39:25]
  assign _T_238 = {_T_233,_T_237}; // @[Cat.scala 29:58]
  assign _T_239 = _T_231[1:0]; // @[LZD.scala 44:32]
  assign _T_240 = _T_239 != 2'h0; // @[LZD.scala 39:14]
  assign _T_241 = _T_239[1]; // @[LZD.scala 39:21]
  assign _T_242 = _T_239[0]; // @[LZD.scala 39:30]
  assign _T_243 = ~ _T_242; // @[LZD.scala 39:27]
  assign _T_244 = _T_241 | _T_243; // @[LZD.scala 39:25]
  assign _T_245 = {_T_240,_T_244}; // @[Cat.scala 29:58]
  assign _T_246 = _T_238[1]; // @[Shift.scala 12:21]
  assign _T_247 = _T_245[1]; // @[Shift.scala 12:21]
  assign _T_248 = _T_246 | _T_247; // @[LZD.scala 49:16]
  assign _T_249 = ~ _T_247; // @[LZD.scala 49:27]
  assign _T_250 = _T_246 | _T_249; // @[LZD.scala 49:25]
  assign _T_251 = _T_238[0:0]; // @[LZD.scala 49:47]
  assign _T_252 = _T_245[0:0]; // @[LZD.scala 49:59]
  assign _T_253 = _T_246 ? _T_251 : _T_252; // @[LZD.scala 49:35]
  assign _T_255 = {_T_248,_T_250,_T_253}; // @[Cat.scala 29:58]
  assign _T_256 = _T_230[1:0]; // @[LZD.scala 44:32]
  assign _T_257 = _T_256 != 2'h0; // @[LZD.scala 39:14]
  assign _T_258 = _T_256[1]; // @[LZD.scala 39:21]
  assign _T_259 = _T_256[0]; // @[LZD.scala 39:30]
  assign _T_260 = ~ _T_259; // @[LZD.scala 39:27]
  assign _T_261 = _T_258 | _T_260; // @[LZD.scala 39:25]
  assign _T_262 = {_T_257,_T_261}; // @[Cat.scala 29:58]
  assign _T_263 = _T_255[2]; // @[Shift.scala 12:21]
  assign _T_265 = _T_255[1:0]; // @[LZD.scala 55:32]
  assign _T_266 = _T_263 ? _T_265 : _T_262; // @[LZD.scala 55:20]
  assign _T_267 = {_T_263,_T_266}; // @[Cat.scala 29:58]
  assign _T_268 = _T_229[3]; // @[Shift.scala 12:21]
  assign _T_270 = _T_229[2:0]; // @[LZD.scala 55:32]
  assign _T_271 = _T_268 ? _T_270 : _T_267; // @[LZD.scala 55:20]
  assign _T_272 = {_T_268,_T_271}; // @[Cat.scala 29:58]
  assign _T_273 = ~ _T_272; // @[convert.scala 21:22]
  assign _T_274 = io_B[12:0]; // @[convert.scala 22:36]
  assign _T_275 = _T_273 < 4'hd; // @[Shift.scala 16:24]
  assign _T_277 = _T_273[3]; // @[Shift.scala 12:21]
  assign _T_278 = _T_274[4:0]; // @[Shift.scala 64:52]
  assign _T_280 = {_T_278,8'h0}; // @[Cat.scala 29:58]
  assign _T_281 = _T_277 ? _T_280 : _T_274; // @[Shift.scala 64:27]
  assign _T_282 = _T_273[2:0]; // @[Shift.scala 66:70]
  assign _T_283 = _T_282[2]; // @[Shift.scala 12:21]
  assign _T_284 = _T_281[8:0]; // @[Shift.scala 64:52]
  assign _T_286 = {_T_284,4'h0}; // @[Cat.scala 29:58]
  assign _T_287 = _T_283 ? _T_286 : _T_281; // @[Shift.scala 64:27]
  assign _T_288 = _T_282[1:0]; // @[Shift.scala 66:70]
  assign _T_289 = _T_288[1]; // @[Shift.scala 12:21]
  assign _T_290 = _T_287[10:0]; // @[Shift.scala 64:52]
  assign _T_292 = {_T_290,2'h0}; // @[Cat.scala 29:58]
  assign _T_293 = _T_289 ? _T_292 : _T_287; // @[Shift.scala 64:27]
  assign _T_294 = _T_288[0:0]; // @[Shift.scala 66:70]
  assign _T_296 = _T_293[11:0]; // @[Shift.scala 64:52]
  assign _T_297 = {_T_296,1'h0}; // @[Cat.scala 29:58]
  assign _T_298 = _T_294 ? _T_297 : _T_293; // @[Shift.scala 64:27]
  assign _T_299 = _T_275 ? _T_298 : 13'h0; // @[Shift.scala 16:10]
  assign _T_300 = _T_299[12:9]; // @[convert.scala 23:34]
  assign decB_fraction = _T_299[8:0]; // @[convert.scala 24:34]
  assign _T_302 = _T_165 == 1'h0; // @[convert.scala 25:26]
  assign _T_304 = _T_165 ? _T_273 : _T_272; // @[convert.scala 25:42]
  assign _T_307 = ~ _T_300; // @[convert.scala 26:67]
  assign _T_308 = _T_163 ? _T_307 : _T_300; // @[convert.scala 26:51]
  assign _T_309 = {_T_302,_T_304,_T_308}; // @[Cat.scala 29:58]
  assign _T_311 = io_B[14:0]; // @[convert.scala 29:56]
  assign _T_312 = _T_311 != 15'h0; // @[convert.scala 29:60]
  assign _T_313 = ~ _T_312; // @[convert.scala 29:41]
  assign decB_isNaR = _T_163 & _T_313; // @[convert.scala 29:39]
  assign _T_316 = _T_163 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_316 & _T_313; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_309); // @[convert.scala 32:24]
  assign _T_324 = ~ _T_1; // @[PositMultiplier.scala 43:34]
  assign _T_326 = {_T_1,_T_324,decA_fraction}; // @[Cat.scala 29:58]
  assign sigA = $signed(_T_326); // @[PositMultiplier.scala 43:61]
  assign _T_327 = ~ _T_163; // @[PositMultiplier.scala 44:34]
  assign _T_329 = {_T_163,_T_327,decB_fraction}; // @[Cat.scala 29:58]
  assign sigB = $signed(_T_329); // @[PositMultiplier.scala 44:61]
  assign _T_330 = $signed(sigA) * $signed(sigB); // @[PositMultiplier.scala 45:25]
  assign sigP = $unsigned(_T_330); // @[PositMultiplier.scala 45:33]
  assign head2 = sigP[21:20]; // @[PositMultiplier.scala 46:28]
  assign _T_331 = head2[1]; // @[PositMultiplier.scala 47:31]
  assign _T_332 = ~ _T_331; // @[PositMultiplier.scala 47:25]
  assign _T_333 = head2[0]; // @[PositMultiplier.scala 47:42]
  assign addTwo = _T_332 & _T_333; // @[PositMultiplier.scala 47:35]
  assign _T_334 = sigP[21]; // @[PositMultiplier.scala 49:23]
  assign _T_335 = sigP[19]; // @[PositMultiplier.scala 49:49]
  assign addOne = _T_334 ^ _T_335; // @[PositMultiplier.scala 49:43]
  assign _T_336 = {addTwo,addOne}; // @[Cat.scala 29:58]
  assign expBias = {1'b0,$signed(_T_336)}; // @[PositMultiplier.scala 50:39]
  assign _T_337 = sigP[18:0]; // @[PositMultiplier.scala 53:81]
  assign _T_338 = sigP[17:0]; // @[PositMultiplier.scala 54:81]
  assign _T_339 = {_T_338, 1'h0}; // @[PositMultiplier.scala 54:104]
  assign frac = addOne ? _T_337 : _T_339; // @[PositMultiplier.scala 51:22]
  assign _T_340 = $signed(decA_scale) + $signed(decB_scale); // @[PositMultiplier.scala 56:30]
  assign _GEN_0 = {{7{expBias[2]}},expBias}; // @[PositMultiplier.scala 56:44]
  assign _T_342 = $signed(_T_340) + $signed(_GEN_0); // @[PositMultiplier.scala 56:44]
  assign mulScale = $signed(_T_342); // @[PositMultiplier.scala 56:44]
  assign underflow = $signed(mulScale) < $signed(-10'she0); // @[PositMultiplier.scala 57:28]
  assign overflow = $signed(mulScale) > $signed(10'she0); // @[PositMultiplier.scala 58:28]
  assign decM_sign = sigP[21:21]; // @[PositMultiplier.scala 62:29]
  assign _T_345 = underflow ? $signed(-10'she0) : $signed(mulScale); // @[Mux.scala 87:16]
  assign _T_346 = overflow ? $signed(10'she0) : $signed(_T_345); // @[Mux.scala 87:16]
  assign decM_fraction = frac[18:10]; // @[PositMultiplier.scala 70:29]
  assign decM_isNaR = decA_isNaR | decB_isNaR; // @[PositMultiplier.scala 71:31]
  assign decM_isZero = decA_isZero | decB_isZero; // @[PositMultiplier.scala 72:32]
  assign grsTmp = frac[9:0]; // @[PositMultiplier.scala 75:30]
  assign _T_350 = grsTmp[9:8]; // @[PositMultiplier.scala 78:32]
  assign _T_351 = grsTmp[7:0]; // @[PositMultiplier.scala 78:48]
  assign _T_352 = _T_351 != 8'h0; // @[PositMultiplier.scala 78:52]
  assign _GEN_1 = _T_346[8:0]; // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  assign decM_scale = $signed(_GEN_1); // @[PositMultiplier.scala 60:23 PositMultiplier.scala 63:17]
  assign _T_355 = decM_scale[3:0]; // @[convert.scala 46:61]
  assign _T_356 = ~ _T_355; // @[convert.scala 46:52]
  assign _T_358 = decM_sign ? _T_356 : _T_355; // @[convert.scala 46:42]
  assign _T_359 = decM_scale[8:4]; // @[convert.scala 48:34]
  assign _T_360 = _T_359[4:4]; // @[convert.scala 49:36]
  assign _T_362 = ~ _T_359; // @[convert.scala 50:36]
  assign _T_363 = $signed(_T_362); // @[convert.scala 50:36]
  assign _T_364 = _T_360 ? $signed(_T_363) : $signed(_T_359); // @[convert.scala 50:28]
  assign _T_365 = _T_360 ^ decM_sign; // @[convert.scala 51:31]
  assign _T_366 = ~ _T_365; // @[convert.scala 52:43]
  assign _T_370 = {_T_366,_T_365,_T_358,decM_fraction,_T_350,_T_352}; // @[Cat.scala 29:58]
  assign _T_371 = $unsigned(_T_364); // @[Shift.scala 39:17]
  assign _T_372 = _T_371 < 5'h12; // @[Shift.scala 39:24]
  assign _T_374 = _T_370[17:16]; // @[Shift.scala 90:30]
  assign _T_375 = _T_370[15:0]; // @[Shift.scala 90:48]
  assign _T_376 = _T_375 != 16'h0; // @[Shift.scala 90:57]
  assign _GEN_2 = {{1'd0}, _T_376}; // @[Shift.scala 90:39]
  assign _T_377 = _T_374 | _GEN_2; // @[Shift.scala 90:39]
  assign _T_378 = _T_371[4]; // @[Shift.scala 12:21]
  assign _T_379 = _T_370[17]; // @[Shift.scala 12:21]
  assign _T_381 = _T_379 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_382 = {_T_381,_T_377}; // @[Cat.scala 29:58]
  assign _T_383 = _T_378 ? _T_382 : _T_370; // @[Shift.scala 91:22]
  assign _T_384 = _T_371[3:0]; // @[Shift.scala 92:77]
  assign _T_385 = _T_383[17:8]; // @[Shift.scala 90:30]
  assign _T_386 = _T_383[7:0]; // @[Shift.scala 90:48]
  assign _T_387 = _T_386 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_3 = {{9'd0}, _T_387}; // @[Shift.scala 90:39]
  assign _T_388 = _T_385 | _GEN_3; // @[Shift.scala 90:39]
  assign _T_389 = _T_384[3]; // @[Shift.scala 12:21]
  assign _T_390 = _T_383[17]; // @[Shift.scala 12:21]
  assign _T_392 = _T_390 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_393 = {_T_392,_T_388}; // @[Cat.scala 29:58]
  assign _T_394 = _T_389 ? _T_393 : _T_383; // @[Shift.scala 91:22]
  assign _T_395 = _T_384[2:0]; // @[Shift.scala 92:77]
  assign _T_396 = _T_394[17:4]; // @[Shift.scala 90:30]
  assign _T_397 = _T_394[3:0]; // @[Shift.scala 90:48]
  assign _T_398 = _T_397 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_4 = {{13'd0}, _T_398}; // @[Shift.scala 90:39]
  assign _T_399 = _T_396 | _GEN_4; // @[Shift.scala 90:39]
  assign _T_400 = _T_395[2]; // @[Shift.scala 12:21]
  assign _T_401 = _T_394[17]; // @[Shift.scala 12:21]
  assign _T_403 = _T_401 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_404 = {_T_403,_T_399}; // @[Cat.scala 29:58]
  assign _T_405 = _T_400 ? _T_404 : _T_394; // @[Shift.scala 91:22]
  assign _T_406 = _T_395[1:0]; // @[Shift.scala 92:77]
  assign _T_407 = _T_405[17:2]; // @[Shift.scala 90:30]
  assign _T_408 = _T_405[1:0]; // @[Shift.scala 90:48]
  assign _T_409 = _T_408 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_5 = {{15'd0}, _T_409}; // @[Shift.scala 90:39]
  assign _T_410 = _T_407 | _GEN_5; // @[Shift.scala 90:39]
  assign _T_411 = _T_406[1]; // @[Shift.scala 12:21]
  assign _T_412 = _T_405[17]; // @[Shift.scala 12:21]
  assign _T_414 = _T_412 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_415 = {_T_414,_T_410}; // @[Cat.scala 29:58]
  assign _T_416 = _T_411 ? _T_415 : _T_405; // @[Shift.scala 91:22]
  assign _T_417 = _T_406[0:0]; // @[Shift.scala 92:77]
  assign _T_418 = _T_416[17:1]; // @[Shift.scala 90:30]
  assign _T_419 = _T_416[0:0]; // @[Shift.scala 90:48]
  assign _GEN_6 = {{16'd0}, _T_419}; // @[Shift.scala 90:39]
  assign _T_421 = _T_418 | _GEN_6; // @[Shift.scala 90:39]
  assign _T_423 = _T_416[17]; // @[Shift.scala 12:21]
  assign _T_424 = {_T_423,_T_421}; // @[Cat.scala 29:58]
  assign _T_425 = _T_417 ? _T_424 : _T_416; // @[Shift.scala 91:22]
  assign _T_428 = _T_379 ? 18'h3ffff : 18'h0; // @[Bitwise.scala 71:12]
  assign _T_429 = _T_372 ? _T_425 : _T_428; // @[Shift.scala 39:10]
  assign _T_430 = _T_429[3]; // @[convert.scala 55:31]
  assign _T_431 = _T_429[2]; // @[convert.scala 56:31]
  assign _T_432 = _T_429[1]; // @[convert.scala 57:31]
  assign _T_433 = _T_429[0]; // @[convert.scala 58:31]
  assign _T_434 = _T_429[17:3]; // @[convert.scala 59:69]
  assign _T_435 = _T_434 != 15'h0; // @[convert.scala 59:81]
  assign _T_436 = ~ _T_435; // @[convert.scala 59:50]
  assign _T_438 = _T_434 == 15'h7fff; // @[convert.scala 60:81]
  assign _T_439 = _T_430 | _T_432; // @[convert.scala 61:44]
  assign _T_440 = _T_439 | _T_433; // @[convert.scala 61:52]
  assign _T_441 = _T_431 & _T_440; // @[convert.scala 61:36]
  assign _T_442 = ~ _T_438; // @[convert.scala 62:63]
  assign _T_443 = _T_442 & _T_441; // @[convert.scala 62:103]
  assign _T_444 = _T_436 | _T_443; // @[convert.scala 62:60]
  assign _GEN_7 = {{14'd0}, _T_444}; // @[convert.scala 63:56]
  assign _T_447 = _T_434 + _GEN_7; // @[convert.scala 63:56]
  assign _T_448 = {decM_sign,_T_447}; // @[Cat.scala 29:58]
  assign _T_450 = decM_isZero ? 16'h0 : _T_448; // @[Mux.scala 87:16]
  assign io_M = decM_isNaR ? 16'h8000 : _T_450; // @[PositMultiplier.scala 86:8]
endmodule
