module PositDivSqrter14_1(
  input         clock,
  input         reset,
  output        io_inReady,
  input         io_inValid,
  input         io_sqrtOp,
  input  [13:0] io_A,
  input  [13:0] io_B,
  output        io_diviValid,
  output        io_sqrtValid,
  output        io_invalidExc,
  output [13:0] io_Q
);
  reg [3:0] cycleNum; // @[PositDivisionSqrt.scala 63:26]
  reg [31:0] _RAND_0;
  reg  sqrtOp_Z; // @[PositDivisionSqrt.scala 65:22]
  reg [31:0] _RAND_1;
  reg  isNaR_Z; // @[PositDivisionSqrt.scala 66:22]
  reg [31:0] _RAND_2;
  reg  isZero_Z; // @[PositDivisionSqrt.scala 67:22]
  reg [31:0] _RAND_3;
  reg [6:0] scale_Z; // @[PositDivisionSqrt.scala 68:22]
  reg [31:0] _RAND_4;
  reg  signB_Z; // @[PositDivisionSqrt.scala 69:28]
  reg [31:0] _RAND_5;
  reg [9:0] fractB_Z; // @[PositDivisionSqrt.scala 70:22]
  reg [31:0] _RAND_6;
  reg [13:0] rem_Z; // @[PositDivisionSqrt.scala 71:22]
  reg [31:0] _RAND_7;
  reg [13:0] sigX_Z; // @[PositDivisionSqrt.scala 72:22]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[convert.scala 18:24]
  wire  _T_2; // @[convert.scala 18:40]
  wire  _T_3; // @[convert.scala 18:36]
  wire [11:0] _T_4; // @[convert.scala 19:24]
  wire [11:0] _T_5; // @[convert.scala 19:43]
  wire [11:0] _T_6; // @[convert.scala 19:39]
  wire [7:0] _T_7; // @[LZD.scala 43:32]
  wire [3:0] _T_8; // @[LZD.scala 43:32]
  wire [1:0] _T_9; // @[LZD.scala 43:32]
  wire  _T_10; // @[LZD.scala 39:14]
  wire  _T_11; // @[LZD.scala 39:21]
  wire  _T_12; // @[LZD.scala 39:30]
  wire  _T_13; // @[LZD.scala 39:27]
  wire  _T_14; // @[LZD.scala 39:25]
  wire [1:0] _T_15; // @[Cat.scala 29:58]
  wire [1:0] _T_16; // @[LZD.scala 44:32]
  wire  _T_17; // @[LZD.scala 39:14]
  wire  _T_18; // @[LZD.scala 39:21]
  wire  _T_19; // @[LZD.scala 39:30]
  wire  _T_20; // @[LZD.scala 39:27]
  wire  _T_21; // @[LZD.scala 39:25]
  wire [1:0] _T_22; // @[Cat.scala 29:58]
  wire  _T_23; // @[Shift.scala 12:21]
  wire  _T_24; // @[Shift.scala 12:21]
  wire  _T_25; // @[LZD.scala 49:16]
  wire  _T_26; // @[LZD.scala 49:27]
  wire  _T_27; // @[LZD.scala 49:25]
  wire  _T_28; // @[LZD.scala 49:47]
  wire  _T_29; // @[LZD.scala 49:59]
  wire  _T_30; // @[LZD.scala 49:35]
  wire [2:0] _T_32; // @[Cat.scala 29:58]
  wire [3:0] _T_33; // @[LZD.scala 44:32]
  wire [1:0] _T_34; // @[LZD.scala 43:32]
  wire  _T_35; // @[LZD.scala 39:14]
  wire  _T_36; // @[LZD.scala 39:21]
  wire  _T_37; // @[LZD.scala 39:30]
  wire  _T_38; // @[LZD.scala 39:27]
  wire  _T_39; // @[LZD.scala 39:25]
  wire [1:0] _T_40; // @[Cat.scala 29:58]
  wire [1:0] _T_41; // @[LZD.scala 44:32]
  wire  _T_42; // @[LZD.scala 39:14]
  wire  _T_43; // @[LZD.scala 39:21]
  wire  _T_44; // @[LZD.scala 39:30]
  wire  _T_45; // @[LZD.scala 39:27]
  wire  _T_46; // @[LZD.scala 39:25]
  wire [1:0] _T_47; // @[Cat.scala 29:58]
  wire  _T_48; // @[Shift.scala 12:21]
  wire  _T_49; // @[Shift.scala 12:21]
  wire  _T_50; // @[LZD.scala 49:16]
  wire  _T_51; // @[LZD.scala 49:27]
  wire  _T_52; // @[LZD.scala 49:25]
  wire  _T_53; // @[LZD.scala 49:47]
  wire  _T_54; // @[LZD.scala 49:59]
  wire  _T_55; // @[LZD.scala 49:35]
  wire [2:0] _T_57; // @[Cat.scala 29:58]
  wire  _T_58; // @[Shift.scala 12:21]
  wire  _T_59; // @[Shift.scala 12:21]
  wire  _T_60; // @[LZD.scala 49:16]
  wire  _T_61; // @[LZD.scala 49:27]
  wire  _T_62; // @[LZD.scala 49:25]
  wire [1:0] _T_63; // @[LZD.scala 49:47]
  wire [1:0] _T_64; // @[LZD.scala 49:59]
  wire [1:0] _T_65; // @[LZD.scala 49:35]
  wire [3:0] _T_67; // @[Cat.scala 29:58]
  wire [3:0] _T_68; // @[LZD.scala 44:32]
  wire [1:0] _T_69; // @[LZD.scala 43:32]
  wire  _T_70; // @[LZD.scala 39:14]
  wire  _T_71; // @[LZD.scala 39:21]
  wire  _T_72; // @[LZD.scala 39:30]
  wire  _T_73; // @[LZD.scala 39:27]
  wire  _T_74; // @[LZD.scala 39:25]
  wire [1:0] _T_75; // @[Cat.scala 29:58]
  wire [1:0] _T_76; // @[LZD.scala 44:32]
  wire  _T_77; // @[LZD.scala 39:14]
  wire  _T_78; // @[LZD.scala 39:21]
  wire  _T_79; // @[LZD.scala 39:30]
  wire  _T_80; // @[LZD.scala 39:27]
  wire  _T_81; // @[LZD.scala 39:25]
  wire [1:0] _T_82; // @[Cat.scala 29:58]
  wire  _T_83; // @[Shift.scala 12:21]
  wire  _T_84; // @[Shift.scala 12:21]
  wire  _T_85; // @[LZD.scala 49:16]
  wire  _T_86; // @[LZD.scala 49:27]
  wire  _T_87; // @[LZD.scala 49:25]
  wire  _T_88; // @[LZD.scala 49:47]
  wire  _T_89; // @[LZD.scala 49:59]
  wire  _T_90; // @[LZD.scala 49:35]
  wire [2:0] _T_92; // @[Cat.scala 29:58]
  wire  _T_93; // @[Shift.scala 12:21]
  wire [2:0] _T_95; // @[LZD.scala 55:32]
  wire [2:0] _T_96; // @[LZD.scala 55:20]
  wire [3:0] _T_97; // @[Cat.scala 29:58]
  wire [3:0] _T_98; // @[convert.scala 21:22]
  wire [10:0] _T_99; // @[convert.scala 22:36]
  wire  _T_100; // @[Shift.scala 16:24]
  wire  _T_102; // @[Shift.scala 12:21]
  wire [2:0] _T_103; // @[Shift.scala 64:52]
  wire [10:0] _T_105; // @[Cat.scala 29:58]
  wire [10:0] _T_106; // @[Shift.scala 64:27]
  wire [2:0] _T_107; // @[Shift.scala 66:70]
  wire  _T_108; // @[Shift.scala 12:21]
  wire [6:0] _T_109; // @[Shift.scala 64:52]
  wire [10:0] _T_111; // @[Cat.scala 29:58]
  wire [10:0] _T_112; // @[Shift.scala 64:27]
  wire [1:0] _T_113; // @[Shift.scala 66:70]
  wire  _T_114; // @[Shift.scala 12:21]
  wire [8:0] _T_115; // @[Shift.scala 64:52]
  wire [10:0] _T_117; // @[Cat.scala 29:58]
  wire [10:0] _T_118; // @[Shift.scala 64:27]
  wire  _T_119; // @[Shift.scala 66:70]
  wire [9:0] _T_121; // @[Shift.scala 64:52]
  wire [10:0] _T_122; // @[Cat.scala 29:58]
  wire [10:0] _T_123; // @[Shift.scala 64:27]
  wire [10:0] _T_124; // @[Shift.scala 16:10]
  wire  _T_125; // @[convert.scala 23:34]
  wire [9:0] decA_fraction; // @[convert.scala 24:34]
  wire  _T_127; // @[convert.scala 25:26]
  wire [3:0] _T_129; // @[convert.scala 25:42]
  wire  _T_132; // @[convert.scala 26:67]
  wire  _T_133; // @[convert.scala 26:51]
  wire [5:0] _T_134; // @[Cat.scala 29:58]
  wire [12:0] _T_136; // @[convert.scala 29:56]
  wire  _T_137; // @[convert.scala 29:60]
  wire  _T_138; // @[convert.scala 29:41]
  wire  decA_isNaR; // @[convert.scala 29:39]
  wire  _T_141; // @[convert.scala 30:19]
  wire  decA_isZero; // @[convert.scala 30:41]
  wire [5:0] decA_scale; // @[convert.scala 32:24]
  wire  _T_150; // @[convert.scala 18:24]
  wire  _T_151; // @[convert.scala 18:40]
  wire  _T_152; // @[convert.scala 18:36]
  wire [11:0] _T_153; // @[convert.scala 19:24]
  wire [11:0] _T_154; // @[convert.scala 19:43]
  wire [11:0] _T_155; // @[convert.scala 19:39]
  wire [7:0] _T_156; // @[LZD.scala 43:32]
  wire [3:0] _T_157; // @[LZD.scala 43:32]
  wire [1:0] _T_158; // @[LZD.scala 43:32]
  wire  _T_159; // @[LZD.scala 39:14]
  wire  _T_160; // @[LZD.scala 39:21]
  wire  _T_161; // @[LZD.scala 39:30]
  wire  _T_162; // @[LZD.scala 39:27]
  wire  _T_163; // @[LZD.scala 39:25]
  wire [1:0] _T_164; // @[Cat.scala 29:58]
  wire [1:0] _T_165; // @[LZD.scala 44:32]
  wire  _T_166; // @[LZD.scala 39:14]
  wire  _T_167; // @[LZD.scala 39:21]
  wire  _T_168; // @[LZD.scala 39:30]
  wire  _T_169; // @[LZD.scala 39:27]
  wire  _T_170; // @[LZD.scala 39:25]
  wire [1:0] _T_171; // @[Cat.scala 29:58]
  wire  _T_172; // @[Shift.scala 12:21]
  wire  _T_173; // @[Shift.scala 12:21]
  wire  _T_174; // @[LZD.scala 49:16]
  wire  _T_175; // @[LZD.scala 49:27]
  wire  _T_176; // @[LZD.scala 49:25]
  wire  _T_177; // @[LZD.scala 49:47]
  wire  _T_178; // @[LZD.scala 49:59]
  wire  _T_179; // @[LZD.scala 49:35]
  wire [2:0] _T_181; // @[Cat.scala 29:58]
  wire [3:0] _T_182; // @[LZD.scala 44:32]
  wire [1:0] _T_183; // @[LZD.scala 43:32]
  wire  _T_184; // @[LZD.scala 39:14]
  wire  _T_185; // @[LZD.scala 39:21]
  wire  _T_186; // @[LZD.scala 39:30]
  wire  _T_187; // @[LZD.scala 39:27]
  wire  _T_188; // @[LZD.scala 39:25]
  wire [1:0] _T_189; // @[Cat.scala 29:58]
  wire [1:0] _T_190; // @[LZD.scala 44:32]
  wire  _T_191; // @[LZD.scala 39:14]
  wire  _T_192; // @[LZD.scala 39:21]
  wire  _T_193; // @[LZD.scala 39:30]
  wire  _T_194; // @[LZD.scala 39:27]
  wire  _T_195; // @[LZD.scala 39:25]
  wire [1:0] _T_196; // @[Cat.scala 29:58]
  wire  _T_197; // @[Shift.scala 12:21]
  wire  _T_198; // @[Shift.scala 12:21]
  wire  _T_199; // @[LZD.scala 49:16]
  wire  _T_200; // @[LZD.scala 49:27]
  wire  _T_201; // @[LZD.scala 49:25]
  wire  _T_202; // @[LZD.scala 49:47]
  wire  _T_203; // @[LZD.scala 49:59]
  wire  _T_204; // @[LZD.scala 49:35]
  wire [2:0] _T_206; // @[Cat.scala 29:58]
  wire  _T_207; // @[Shift.scala 12:21]
  wire  _T_208; // @[Shift.scala 12:21]
  wire  _T_209; // @[LZD.scala 49:16]
  wire  _T_210; // @[LZD.scala 49:27]
  wire  _T_211; // @[LZD.scala 49:25]
  wire [1:0] _T_212; // @[LZD.scala 49:47]
  wire [1:0] _T_213; // @[LZD.scala 49:59]
  wire [1:0] _T_214; // @[LZD.scala 49:35]
  wire [3:0] _T_216; // @[Cat.scala 29:58]
  wire [3:0] _T_217; // @[LZD.scala 44:32]
  wire [1:0] _T_218; // @[LZD.scala 43:32]
  wire  _T_219; // @[LZD.scala 39:14]
  wire  _T_220; // @[LZD.scala 39:21]
  wire  _T_221; // @[LZD.scala 39:30]
  wire  _T_222; // @[LZD.scala 39:27]
  wire  _T_223; // @[LZD.scala 39:25]
  wire [1:0] _T_224; // @[Cat.scala 29:58]
  wire [1:0] _T_225; // @[LZD.scala 44:32]
  wire  _T_226; // @[LZD.scala 39:14]
  wire  _T_227; // @[LZD.scala 39:21]
  wire  _T_228; // @[LZD.scala 39:30]
  wire  _T_229; // @[LZD.scala 39:27]
  wire  _T_230; // @[LZD.scala 39:25]
  wire [1:0] _T_231; // @[Cat.scala 29:58]
  wire  _T_232; // @[Shift.scala 12:21]
  wire  _T_233; // @[Shift.scala 12:21]
  wire  _T_234; // @[LZD.scala 49:16]
  wire  _T_235; // @[LZD.scala 49:27]
  wire  _T_236; // @[LZD.scala 49:25]
  wire  _T_237; // @[LZD.scala 49:47]
  wire  _T_238; // @[LZD.scala 49:59]
  wire  _T_239; // @[LZD.scala 49:35]
  wire [2:0] _T_241; // @[Cat.scala 29:58]
  wire  _T_242; // @[Shift.scala 12:21]
  wire [2:0] _T_244; // @[LZD.scala 55:32]
  wire [2:0] _T_245; // @[LZD.scala 55:20]
  wire [3:0] _T_246; // @[Cat.scala 29:58]
  wire [3:0] _T_247; // @[convert.scala 21:22]
  wire [10:0] _T_248; // @[convert.scala 22:36]
  wire  _T_249; // @[Shift.scala 16:24]
  wire  _T_251; // @[Shift.scala 12:21]
  wire [2:0] _T_252; // @[Shift.scala 64:52]
  wire [10:0] _T_254; // @[Cat.scala 29:58]
  wire [10:0] _T_255; // @[Shift.scala 64:27]
  wire [2:0] _T_256; // @[Shift.scala 66:70]
  wire  _T_257; // @[Shift.scala 12:21]
  wire [6:0] _T_258; // @[Shift.scala 64:52]
  wire [10:0] _T_260; // @[Cat.scala 29:58]
  wire [10:0] _T_261; // @[Shift.scala 64:27]
  wire [1:0] _T_262; // @[Shift.scala 66:70]
  wire  _T_263; // @[Shift.scala 12:21]
  wire [8:0] _T_264; // @[Shift.scala 64:52]
  wire [10:0] _T_266; // @[Cat.scala 29:58]
  wire [10:0] _T_267; // @[Shift.scala 64:27]
  wire  _T_268; // @[Shift.scala 66:70]
  wire [9:0] _T_270; // @[Shift.scala 64:52]
  wire [10:0] _T_271; // @[Cat.scala 29:58]
  wire [10:0] _T_272; // @[Shift.scala 64:27]
  wire [10:0] _T_273; // @[Shift.scala 16:10]
  wire  _T_274; // @[convert.scala 23:34]
  wire [9:0] decB_fraction; // @[convert.scala 24:34]
  wire  _T_276; // @[convert.scala 25:26]
  wire [3:0] _T_278; // @[convert.scala 25:42]
  wire  _T_281; // @[convert.scala 26:67]
  wire  _T_282; // @[convert.scala 26:51]
  wire [5:0] _T_283; // @[Cat.scala 29:58]
  wire [12:0] _T_285; // @[convert.scala 29:56]
  wire  _T_286; // @[convert.scala 29:60]
  wire  _T_287; // @[convert.scala 29:41]
  wire  decB_isNaR; // @[convert.scala 29:39]
  wire  _T_290; // @[convert.scala 30:19]
  wire  decB_isZero; // @[convert.scala 30:41]
  wire [5:0] decB_scale; // @[convert.scala 32:24]
  wire [2:0] _T_299; // @[Bitwise.scala 71:12]
  wire  _T_300; // @[PositDivisionSqrt.scala 80:40]
  wire [13:0] sigA_S; // @[Cat.scala 29:58]
  wire  _T_302; // @[PositDivisionSqrt.scala 82:31]
  wire [13:0] sigB_S; // @[Cat.scala 29:58]
  wire  _T_305; // @[PositDivisionSqrt.scala 85:25]
  wire  invalidSqrt; // @[PositDivisionSqrt.scala 85:37]
  wire  _T_306; // @[PositDivisionSqrt.scala 88:42]
  wire  _T_307; // @[PositDivisionSqrt.scala 89:42]
  wire  _T_308; // @[PositDivisionSqrt.scala 89:56]
  wire  _T_309; // @[PositDivisionSqrt.scala 94:46]
  wire  _T_310; // @[PositDivisionSqrt.scala 94:43]
  wire  _T_311; // @[PositDivisionSqrt.scala 94:62]
  wire  _T_312; // @[PositDivisionSqrt.scala 94:59]
  wire  specialCaseA_S; // @[PositDivisionSqrt.scala 97:38]
  wire  specialCaseB_S; // @[PositDivisionSqrt.scala 98:38]
  wire  _T_313; // @[PositDivisionSqrt.scala 99:27]
  wire  _T_314; // @[PositDivisionSqrt.scala 99:46]
  wire  normalCase_S_div; // @[PositDivisionSqrt.scala 99:43]
  wire  normalCase_S_sqrt; // @[PositDivisionSqrt.scala 100:43]
  wire  normalCase_S; // @[PositDivisionSqrt.scala 101:30]
  wire [6:0] sExpQuot_S_div; // @[PositDivisionSqrt.scala 103:38]
  wire  _T_317; // @[PositDivisionSqrt.scala 104:50]
  wire  oddSqrt_S; // @[PositDivisionSqrt.scala 104:37]
  wire  idle; // @[PositDivisionSqrt.scala 109:39]
  wire  ready; // @[PositDivisionSqrt.scala 110:39]
  wire  entering; // @[PositDivisionSqrt.scala 111:35]
  wire  entering_normalCase; // @[PositDivisionSqrt.scala 112:38]
  wire  _T_318; // @[PositDivisionSqrt.scala 113:35]
  wire  _T_319; // @[PositDivisionSqrt.scala 113:58]
  wire  scaleNotChange; // @[PositDivisionSqrt.scala 113:50]
  wire  _T_320; // @[PositDivisionSqrt.scala 114:39]
  wire  skipCycle2; // @[PositDivisionSqrt.scala 114:48]
  wire  _T_321; // @[PositDivisionSqrt.scala 116:8]
  wire  _T_322; // @[PositDivisionSqrt.scala 116:14]
  wire  _T_323; // @[PositDivisionSqrt.scala 117:32]
  wire  _T_324; // @[PositDivisionSqrt.scala 117:30]
  wire [3:0] _T_326; // @[PositDivisionSqrt.scala 119:26]
  wire [3:0] _T_327; // @[PositDivisionSqrt.scala 118:20]
  wire [3:0] _GEN_9; // @[PositDivisionSqrt.scala 117:64]
  wire [3:0] _T_328; // @[PositDivisionSqrt.scala 117:64]
  wire  _T_330; // @[PositDivisionSqrt.scala 123:30]
  wire  _T_331; // @[PositDivisionSqrt.scala 123:27]
  wire [3:0] _T_333; // @[PositDivisionSqrt.scala 123:52]
  wire [3:0] _T_334; // @[PositDivisionSqrt.scala 123:20]
  wire [3:0] _T_335; // @[PositDivisionSqrt.scala 122:64]
  wire  _T_337; // @[PositDivisionSqrt.scala 124:27]
  wire [3:0] _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  wire [3:0] _T_339; // @[PositDivisionSqrt.scala 123:64]
  wire [4:0] _T_340; // @[PositDivisionSqrt.scala 134:42]
  wire  _T_342; // @[PositDivisionSqrt.scala 137:31]
  wire  _T_343; // @[PositDivisionSqrt.scala 137:28]
  wire [15:0] _T_344; // @[PositDivisionSqrt.scala 146:22]
  wire [13:0] _T_345; // @[PositDivisionSqrt.scala 146:35]
  wire  _T_346; // @[PositDivisionSqrt.scala 148:26]
  wire  _T_347; // @[PositDivisionSqrt.scala 148:23]
  wire [13:0] _T_348; // @[PositDivisionSqrt.scala 148:16]
  wire  _T_349; // @[PositDivisionSqrt.scala 149:23]
  wire [14:0] _T_350; // @[PositDivisionSqrt.scala 149:46]
  wire [13:0] _T_351; // @[PositDivisionSqrt.scala 149:56]
  wire [13:0] _T_352; // @[PositDivisionSqrt.scala 149:16]
  wire [13:0] _T_353; // @[PositDivisionSqrt.scala 148:66]
  wire  _T_354; // @[PositDivisionSqrt.scala 150:17]
  wire [13:0] _T_355; // @[PositDivisionSqrt.scala 150:16]
  wire [13:0] rem; // @[PositDivisionSqrt.scala 149:66]
  wire  _T_357; // @[PositDivisionSqrt.scala 152:29]
  wire [13:0] _T_358; // @[PositDivisionSqrt.scala 152:22]
  wire  _T_359; // @[PositDivisionSqrt.scala 153:29]
  wire [10:0] _T_360; // @[PositDivisionSqrt.scala 153:22]
  wire [13:0] _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  wire [13:0] _T_361; // @[PositDivisionSqrt.scala 152:93]
  wire  _T_363; // @[PositDivisionSqrt.scala 154:33]
  wire  _T_364; // @[PositDivisionSqrt.scala 154:30]
  wire  _T_365; // @[PositDivisionSqrt.scala 154:57]
  wire [13:0] _T_368; // @[Cat.scala 29:58]
  wire [13:0] _T_369; // @[PositDivisionSqrt.scala 154:22]
  wire [13:0] _T_370; // @[PositDivisionSqrt.scala 153:93]
  wire  _T_372; // @[PositDivisionSqrt.scala 155:30]
  wire  _T_373; // @[PositDivisionSqrt.scala 156:79]
  wire [9:0] _T_375; // @[Bitwise.scala 71:12]
  wire [12:0] bitMask; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  wire [12:0] _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  wire [12:0] _T_376; // @[PositDivisionSqrt.scala 156:53]
  wire [13:0] _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  wire [13:0] _T_377; // @[PositDivisionSqrt.scala 155:51]
  wire [11:0] _T_378; // @[PositDivisionSqrt.scala 157:53]
  wire [13:0] _GEN_14; // @[PositDivisionSqrt.scala 156:85]
  wire [13:0] _T_379; // @[PositDivisionSqrt.scala 156:85]
  wire [13:0] _T_380; // @[PositDivisionSqrt.scala 155:22]
  wire [13:0] trialTerm; // @[PositDivisionSqrt.scala 154:93]
  wire  _T_382; // @[PositDivisionSqrt.scala 162:56]
  wire  _T_383; // @[PositDivisionSqrt.scala 162:40]
  wire [13:0] _T_386; // @[PositDivisionSqrt.scala 163:97]
  wire [13:0] _T_388; // @[PositDivisionSqrt.scala 164:97]
  wire [13:0] _T_389; // @[PositDivisionSqrt.scala 161:92]
  wire [14:0] _T_394; // @[PositDivisionSqrt.scala 168:98]
  wire [13:0] _T_395; // @[PositDivisionSqrt.scala 168:108]
  wire [13:0] _T_397; // @[PositDivisionSqrt.scala 168:112]
  wire [13:0] _T_401; // @[PositDivisionSqrt.scala 169:112]
  wire [13:0] _T_402; // @[PositDivisionSqrt.scala 166:26]
  wire [13:0] trialRem; // @[PositDivisionSqrt.scala 159:27]
  wire  _T_403; // @[PositDivisionSqrt.scala 173:35]
  wire  trIsZero; // @[PositDivisionSqrt.scala 173:25]
  wire  _T_404; // @[PositDivisionSqrt.scala 174:30]
  wire  remIsZero; // @[PositDivisionSqrt.scala 174:25]
  wire  _T_406; // @[PositDivisionSqrt.scala 176:64]
  wire  _T_407; // @[PositDivisionSqrt.scala 176:49]
  wire  _T_408; // @[PositDivisionSqrt.scala 176:29]
  wire  _T_409; // @[PositDivisionSqrt.scala 178:61]
  wire  _T_410; // @[PositDivisionSqrt.scala 178:49]
  wire  _T_412; // @[Mux.scala 87:16]
  wire  newBit; // @[Mux.scala 87:16]
  wire  _T_413; // @[PositDivisionSqrt.scala 183:41]
  wire  _T_414; // @[PositDivisionSqrt.scala 183:51]
  wire  _T_415; // @[PositDivisionSqrt.scala 183:48]
  wire  _T_416; // @[PositDivisionSqrt.scala 183:28]
  wire  _T_419; // @[PositDivisionSqrt.scala 187:39]
  wire  _T_420; // @[PositDivisionSqrt.scala 187:28]
  wire [13:0] _T_423; // @[PositDivisionSqrt.scala 188:47]
  wire [13:0] _T_424; // @[PositDivisionSqrt.scala 188:18]
  wire [11:0] _T_426; // @[PositDivisionSqrt.scala 189:18]
  wire [13:0] _GEN_15; // @[PositDivisionSqrt.scala 188:72]
  wire [13:0] _T_427; // @[PositDivisionSqrt.scala 188:72]
  wire [13:0] _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  wire [13:0] _T_429; // @[PositDivisionSqrt.scala 190:47]
  wire [13:0] _T_430; // @[PositDivisionSqrt.scala 190:18]
  wire [13:0] _T_431; // @[PositDivisionSqrt.scala 189:72]
  wire [1:0] _T_433; // @[PositDivisionSqrt.scala 196:53]
  wire [1:0] sigXBias; // @[PositDivisionSqrt.scala 196:21]
  wire [13:0] _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  wire [13:0] realSigX; // @[PositDivisionSqrt.scala 197:25]
  wire [9:0] _T_436; // @[PositDivisionSqrt.scala 200:97]
  wire [9:0] _T_437; // @[PositDivisionSqrt.scala 201:97]
  wire [9:0] realFrac; // @[PositDivisionSqrt.scala 198:21]
  wire  _T_438; // @[PositDivisionSqrt.scala 205:33]
  wire  _T_439; // @[PositDivisionSqrt.scala 205:58]
  wire  _T_440; // @[PositDivisionSqrt.scala 205:48]
  wire  scaleNeedSub; // @[PositDivisionSqrt.scala 205:23]
  wire  _T_442; // @[PositDivisionSqrt.scala 206:56]
  wire  notNeedSubTwo; // @[PositDivisionSqrt.scala 206:46]
  wire  scaleSubOne; // @[PositDivisionSqrt.scala 207:36]
  wire  _T_443; // @[PositDivisionSqrt.scala 208:38]
  wire  scaleSubTwo; // @[PositDivisionSqrt.scala 208:36]
  wire [1:0] _T_444; // @[Cat.scala 29:58]
  wire [2:0] _T_445; // @[PositDivisionSqrt.scala 209:63]
  wire [6:0] _GEN_18; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] _T_447; // @[PositDivisionSqrt.scala 209:31]
  wire [6:0] realExp; // @[PositDivisionSqrt.scala 209:31]
  wire  underflow; // @[PositDivisionSqrt.scala 210:31]
  wire  overflow; // @[PositDivisionSqrt.scala 211:31]
  wire  decQ_sign; // @[PositDivisionSqrt.scala 215:33]
  wire [6:0] _T_449; // @[Mux.scala 87:16]
  wire [6:0] _T_450; // @[Mux.scala 87:16]
  wire  outValid; // @[PositDivisionSqrt.scala 229:28]
  wire [5:0] _GEN_19; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire [5:0] decQ_scale; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  wire  _T_455; // @[convert.scala 46:61]
  wire  _T_456; // @[convert.scala 46:52]
  wire  _T_458; // @[convert.scala 46:42]
  wire [4:0] _T_459; // @[convert.scala 48:34]
  wire  _T_460; // @[convert.scala 49:36]
  wire [4:0] _T_462; // @[convert.scala 50:36]
  wire [4:0] _T_463; // @[convert.scala 50:36]
  wire [4:0] _T_464; // @[convert.scala 50:28]
  wire  _T_465; // @[convert.scala 51:31]
  wire  _T_466; // @[convert.scala 52:43]
  wire [15:0] _T_470; // @[Cat.scala 29:58]
  wire [4:0] _T_471; // @[Shift.scala 39:17]
  wire  _T_472; // @[Shift.scala 39:24]
  wire [3:0] _T_473; // @[Shift.scala 40:44]
  wire [7:0] _T_474; // @[Shift.scala 90:30]
  wire [7:0] _T_475; // @[Shift.scala 90:48]
  wire  _T_476; // @[Shift.scala 90:57]
  wire [7:0] _GEN_20; // @[Shift.scala 90:39]
  wire [7:0] _T_477; // @[Shift.scala 90:39]
  wire  _T_478; // @[Shift.scala 12:21]
  wire  _T_479; // @[Shift.scala 12:21]
  wire [7:0] _T_481; // @[Bitwise.scala 71:12]
  wire [15:0] _T_482; // @[Cat.scala 29:58]
  wire [15:0] _T_483; // @[Shift.scala 91:22]
  wire [2:0] _T_484; // @[Shift.scala 92:77]
  wire [11:0] _T_485; // @[Shift.scala 90:30]
  wire [3:0] _T_486; // @[Shift.scala 90:48]
  wire  _T_487; // @[Shift.scala 90:57]
  wire [11:0] _GEN_21; // @[Shift.scala 90:39]
  wire [11:0] _T_488; // @[Shift.scala 90:39]
  wire  _T_489; // @[Shift.scala 12:21]
  wire  _T_490; // @[Shift.scala 12:21]
  wire [3:0] _T_492; // @[Bitwise.scala 71:12]
  wire [15:0] _T_493; // @[Cat.scala 29:58]
  wire [15:0] _T_494; // @[Shift.scala 91:22]
  wire [1:0] _T_495; // @[Shift.scala 92:77]
  wire [13:0] _T_496; // @[Shift.scala 90:30]
  wire [1:0] _T_497; // @[Shift.scala 90:48]
  wire  _T_498; // @[Shift.scala 90:57]
  wire [13:0] _GEN_22; // @[Shift.scala 90:39]
  wire [13:0] _T_499; // @[Shift.scala 90:39]
  wire  _T_500; // @[Shift.scala 12:21]
  wire  _T_501; // @[Shift.scala 12:21]
  wire [1:0] _T_503; // @[Bitwise.scala 71:12]
  wire [15:0] _T_504; // @[Cat.scala 29:58]
  wire [15:0] _T_505; // @[Shift.scala 91:22]
  wire  _T_506; // @[Shift.scala 92:77]
  wire [14:0] _T_507; // @[Shift.scala 90:30]
  wire  _T_508; // @[Shift.scala 90:48]
  wire [14:0] _GEN_23; // @[Shift.scala 90:39]
  wire [14:0] _T_510; // @[Shift.scala 90:39]
  wire  _T_512; // @[Shift.scala 12:21]
  wire [15:0] _T_513; // @[Cat.scala 29:58]
  wire [15:0] _T_514; // @[Shift.scala 91:22]
  wire [15:0] _T_517; // @[Bitwise.scala 71:12]
  wire [15:0] _T_518; // @[Shift.scala 39:10]
  wire  _T_519; // @[convert.scala 55:31]
  wire  _T_520; // @[convert.scala 56:31]
  wire  _T_521; // @[convert.scala 57:31]
  wire  _T_522; // @[convert.scala 58:31]
  wire [12:0] _T_523; // @[convert.scala 59:69]
  wire  _T_524; // @[convert.scala 59:81]
  wire  _T_525; // @[convert.scala 59:50]
  wire  _T_527; // @[convert.scala 60:81]
  wire  _T_528; // @[convert.scala 61:44]
  wire  _T_529; // @[convert.scala 61:52]
  wire  _T_530; // @[convert.scala 61:36]
  wire  _T_531; // @[convert.scala 62:63]
  wire  _T_532; // @[convert.scala 62:103]
  wire  _T_533; // @[convert.scala 62:60]
  wire [12:0] _GEN_24; // @[convert.scala 63:56]
  wire [12:0] _T_536; // @[convert.scala 63:56]
  wire [13:0] _T_537; // @[Cat.scala 29:58]
  wire [13:0] _T_539; // @[Mux.scala 87:16]
  assign _T_1 = io_A[13]; // @[convert.scala 18:24]
  assign _T_2 = io_A[12]; // @[convert.scala 18:40]
  assign _T_3 = _T_1 ^ _T_2; // @[convert.scala 18:36]
  assign _T_4 = io_A[12:1]; // @[convert.scala 19:24]
  assign _T_5 = io_A[11:0]; // @[convert.scala 19:43]
  assign _T_6 = _T_4 ^ _T_5; // @[convert.scala 19:39]
  assign _T_7 = _T_6[11:4]; // @[LZD.scala 43:32]
  assign _T_8 = _T_7[7:4]; // @[LZD.scala 43:32]
  assign _T_9 = _T_8[3:2]; // @[LZD.scala 43:32]
  assign _T_10 = _T_9 != 2'h0; // @[LZD.scala 39:14]
  assign _T_11 = _T_9[1]; // @[LZD.scala 39:21]
  assign _T_12 = _T_9[0]; // @[LZD.scala 39:30]
  assign _T_13 = ~ _T_12; // @[LZD.scala 39:27]
  assign _T_14 = _T_11 | _T_13; // @[LZD.scala 39:25]
  assign _T_15 = {_T_10,_T_14}; // @[Cat.scala 29:58]
  assign _T_16 = _T_8[1:0]; // @[LZD.scala 44:32]
  assign _T_17 = _T_16 != 2'h0; // @[LZD.scala 39:14]
  assign _T_18 = _T_16[1]; // @[LZD.scala 39:21]
  assign _T_19 = _T_16[0]; // @[LZD.scala 39:30]
  assign _T_20 = ~ _T_19; // @[LZD.scala 39:27]
  assign _T_21 = _T_18 | _T_20; // @[LZD.scala 39:25]
  assign _T_22 = {_T_17,_T_21}; // @[Cat.scala 29:58]
  assign _T_23 = _T_15[1]; // @[Shift.scala 12:21]
  assign _T_24 = _T_22[1]; // @[Shift.scala 12:21]
  assign _T_25 = _T_23 | _T_24; // @[LZD.scala 49:16]
  assign _T_26 = ~ _T_24; // @[LZD.scala 49:27]
  assign _T_27 = _T_23 | _T_26; // @[LZD.scala 49:25]
  assign _T_28 = _T_15[0:0]; // @[LZD.scala 49:47]
  assign _T_29 = _T_22[0:0]; // @[LZD.scala 49:59]
  assign _T_30 = _T_23 ? _T_28 : _T_29; // @[LZD.scala 49:35]
  assign _T_32 = {_T_25,_T_27,_T_30}; // @[Cat.scala 29:58]
  assign _T_33 = _T_7[3:0]; // @[LZD.scala 44:32]
  assign _T_34 = _T_33[3:2]; // @[LZD.scala 43:32]
  assign _T_35 = _T_34 != 2'h0; // @[LZD.scala 39:14]
  assign _T_36 = _T_34[1]; // @[LZD.scala 39:21]
  assign _T_37 = _T_34[0]; // @[LZD.scala 39:30]
  assign _T_38 = ~ _T_37; // @[LZD.scala 39:27]
  assign _T_39 = _T_36 | _T_38; // @[LZD.scala 39:25]
  assign _T_40 = {_T_35,_T_39}; // @[Cat.scala 29:58]
  assign _T_41 = _T_33[1:0]; // @[LZD.scala 44:32]
  assign _T_42 = _T_41 != 2'h0; // @[LZD.scala 39:14]
  assign _T_43 = _T_41[1]; // @[LZD.scala 39:21]
  assign _T_44 = _T_41[0]; // @[LZD.scala 39:30]
  assign _T_45 = ~ _T_44; // @[LZD.scala 39:27]
  assign _T_46 = _T_43 | _T_45; // @[LZD.scala 39:25]
  assign _T_47 = {_T_42,_T_46}; // @[Cat.scala 29:58]
  assign _T_48 = _T_40[1]; // @[Shift.scala 12:21]
  assign _T_49 = _T_47[1]; // @[Shift.scala 12:21]
  assign _T_50 = _T_48 | _T_49; // @[LZD.scala 49:16]
  assign _T_51 = ~ _T_49; // @[LZD.scala 49:27]
  assign _T_52 = _T_48 | _T_51; // @[LZD.scala 49:25]
  assign _T_53 = _T_40[0:0]; // @[LZD.scala 49:47]
  assign _T_54 = _T_47[0:0]; // @[LZD.scala 49:59]
  assign _T_55 = _T_48 ? _T_53 : _T_54; // @[LZD.scala 49:35]
  assign _T_57 = {_T_50,_T_52,_T_55}; // @[Cat.scala 29:58]
  assign _T_58 = _T_32[2]; // @[Shift.scala 12:21]
  assign _T_59 = _T_57[2]; // @[Shift.scala 12:21]
  assign _T_60 = _T_58 | _T_59; // @[LZD.scala 49:16]
  assign _T_61 = ~ _T_59; // @[LZD.scala 49:27]
  assign _T_62 = _T_58 | _T_61; // @[LZD.scala 49:25]
  assign _T_63 = _T_32[1:0]; // @[LZD.scala 49:47]
  assign _T_64 = _T_57[1:0]; // @[LZD.scala 49:59]
  assign _T_65 = _T_58 ? _T_63 : _T_64; // @[LZD.scala 49:35]
  assign _T_67 = {_T_60,_T_62,_T_65}; // @[Cat.scala 29:58]
  assign _T_68 = _T_6[3:0]; // @[LZD.scala 44:32]
  assign _T_69 = _T_68[3:2]; // @[LZD.scala 43:32]
  assign _T_70 = _T_69 != 2'h0; // @[LZD.scala 39:14]
  assign _T_71 = _T_69[1]; // @[LZD.scala 39:21]
  assign _T_72 = _T_69[0]; // @[LZD.scala 39:30]
  assign _T_73 = ~ _T_72; // @[LZD.scala 39:27]
  assign _T_74 = _T_71 | _T_73; // @[LZD.scala 39:25]
  assign _T_75 = {_T_70,_T_74}; // @[Cat.scala 29:58]
  assign _T_76 = _T_68[1:0]; // @[LZD.scala 44:32]
  assign _T_77 = _T_76 != 2'h0; // @[LZD.scala 39:14]
  assign _T_78 = _T_76[1]; // @[LZD.scala 39:21]
  assign _T_79 = _T_76[0]; // @[LZD.scala 39:30]
  assign _T_80 = ~ _T_79; // @[LZD.scala 39:27]
  assign _T_81 = _T_78 | _T_80; // @[LZD.scala 39:25]
  assign _T_82 = {_T_77,_T_81}; // @[Cat.scala 29:58]
  assign _T_83 = _T_75[1]; // @[Shift.scala 12:21]
  assign _T_84 = _T_82[1]; // @[Shift.scala 12:21]
  assign _T_85 = _T_83 | _T_84; // @[LZD.scala 49:16]
  assign _T_86 = ~ _T_84; // @[LZD.scala 49:27]
  assign _T_87 = _T_83 | _T_86; // @[LZD.scala 49:25]
  assign _T_88 = _T_75[0:0]; // @[LZD.scala 49:47]
  assign _T_89 = _T_82[0:0]; // @[LZD.scala 49:59]
  assign _T_90 = _T_83 ? _T_88 : _T_89; // @[LZD.scala 49:35]
  assign _T_92 = {_T_85,_T_87,_T_90}; // @[Cat.scala 29:58]
  assign _T_93 = _T_67[3]; // @[Shift.scala 12:21]
  assign _T_95 = _T_67[2:0]; // @[LZD.scala 55:32]
  assign _T_96 = _T_93 ? _T_95 : _T_92; // @[LZD.scala 55:20]
  assign _T_97 = {_T_93,_T_96}; // @[Cat.scala 29:58]
  assign _T_98 = ~ _T_97; // @[convert.scala 21:22]
  assign _T_99 = io_A[10:0]; // @[convert.scala 22:36]
  assign _T_100 = _T_98 < 4'hb; // @[Shift.scala 16:24]
  assign _T_102 = _T_98[3]; // @[Shift.scala 12:21]
  assign _T_103 = _T_99[2:0]; // @[Shift.scala 64:52]
  assign _T_105 = {_T_103,8'h0}; // @[Cat.scala 29:58]
  assign _T_106 = _T_102 ? _T_105 : _T_99; // @[Shift.scala 64:27]
  assign _T_107 = _T_98[2:0]; // @[Shift.scala 66:70]
  assign _T_108 = _T_107[2]; // @[Shift.scala 12:21]
  assign _T_109 = _T_106[6:0]; // @[Shift.scala 64:52]
  assign _T_111 = {_T_109,4'h0}; // @[Cat.scala 29:58]
  assign _T_112 = _T_108 ? _T_111 : _T_106; // @[Shift.scala 64:27]
  assign _T_113 = _T_107[1:0]; // @[Shift.scala 66:70]
  assign _T_114 = _T_113[1]; // @[Shift.scala 12:21]
  assign _T_115 = _T_112[8:0]; // @[Shift.scala 64:52]
  assign _T_117 = {_T_115,2'h0}; // @[Cat.scala 29:58]
  assign _T_118 = _T_114 ? _T_117 : _T_112; // @[Shift.scala 64:27]
  assign _T_119 = _T_113[0:0]; // @[Shift.scala 66:70]
  assign _T_121 = _T_118[9:0]; // @[Shift.scala 64:52]
  assign _T_122 = {_T_121,1'h0}; // @[Cat.scala 29:58]
  assign _T_123 = _T_119 ? _T_122 : _T_118; // @[Shift.scala 64:27]
  assign _T_124 = _T_100 ? _T_123 : 11'h0; // @[Shift.scala 16:10]
  assign _T_125 = _T_124[10:10]; // @[convert.scala 23:34]
  assign decA_fraction = _T_124[9:0]; // @[convert.scala 24:34]
  assign _T_127 = _T_3 == 1'h0; // @[convert.scala 25:26]
  assign _T_129 = _T_3 ? _T_98 : _T_97; // @[convert.scala 25:42]
  assign _T_132 = ~ _T_125; // @[convert.scala 26:67]
  assign _T_133 = _T_1 ? _T_132 : _T_125; // @[convert.scala 26:51]
  assign _T_134 = {_T_127,_T_129,_T_133}; // @[Cat.scala 29:58]
  assign _T_136 = io_A[12:0]; // @[convert.scala 29:56]
  assign _T_137 = _T_136 != 13'h0; // @[convert.scala 29:60]
  assign _T_138 = ~ _T_137; // @[convert.scala 29:41]
  assign decA_isNaR = _T_1 & _T_138; // @[convert.scala 29:39]
  assign _T_141 = _T_1 == 1'h0; // @[convert.scala 30:19]
  assign decA_isZero = _T_141 & _T_138; // @[convert.scala 30:41]
  assign decA_scale = $signed(_T_134); // @[convert.scala 32:24]
  assign _T_150 = io_B[13]; // @[convert.scala 18:24]
  assign _T_151 = io_B[12]; // @[convert.scala 18:40]
  assign _T_152 = _T_150 ^ _T_151; // @[convert.scala 18:36]
  assign _T_153 = io_B[12:1]; // @[convert.scala 19:24]
  assign _T_154 = io_B[11:0]; // @[convert.scala 19:43]
  assign _T_155 = _T_153 ^ _T_154; // @[convert.scala 19:39]
  assign _T_156 = _T_155[11:4]; // @[LZD.scala 43:32]
  assign _T_157 = _T_156[7:4]; // @[LZD.scala 43:32]
  assign _T_158 = _T_157[3:2]; // @[LZD.scala 43:32]
  assign _T_159 = _T_158 != 2'h0; // @[LZD.scala 39:14]
  assign _T_160 = _T_158[1]; // @[LZD.scala 39:21]
  assign _T_161 = _T_158[0]; // @[LZD.scala 39:30]
  assign _T_162 = ~ _T_161; // @[LZD.scala 39:27]
  assign _T_163 = _T_160 | _T_162; // @[LZD.scala 39:25]
  assign _T_164 = {_T_159,_T_163}; // @[Cat.scala 29:58]
  assign _T_165 = _T_157[1:0]; // @[LZD.scala 44:32]
  assign _T_166 = _T_165 != 2'h0; // @[LZD.scala 39:14]
  assign _T_167 = _T_165[1]; // @[LZD.scala 39:21]
  assign _T_168 = _T_165[0]; // @[LZD.scala 39:30]
  assign _T_169 = ~ _T_168; // @[LZD.scala 39:27]
  assign _T_170 = _T_167 | _T_169; // @[LZD.scala 39:25]
  assign _T_171 = {_T_166,_T_170}; // @[Cat.scala 29:58]
  assign _T_172 = _T_164[1]; // @[Shift.scala 12:21]
  assign _T_173 = _T_171[1]; // @[Shift.scala 12:21]
  assign _T_174 = _T_172 | _T_173; // @[LZD.scala 49:16]
  assign _T_175 = ~ _T_173; // @[LZD.scala 49:27]
  assign _T_176 = _T_172 | _T_175; // @[LZD.scala 49:25]
  assign _T_177 = _T_164[0:0]; // @[LZD.scala 49:47]
  assign _T_178 = _T_171[0:0]; // @[LZD.scala 49:59]
  assign _T_179 = _T_172 ? _T_177 : _T_178; // @[LZD.scala 49:35]
  assign _T_181 = {_T_174,_T_176,_T_179}; // @[Cat.scala 29:58]
  assign _T_182 = _T_156[3:0]; // @[LZD.scala 44:32]
  assign _T_183 = _T_182[3:2]; // @[LZD.scala 43:32]
  assign _T_184 = _T_183 != 2'h0; // @[LZD.scala 39:14]
  assign _T_185 = _T_183[1]; // @[LZD.scala 39:21]
  assign _T_186 = _T_183[0]; // @[LZD.scala 39:30]
  assign _T_187 = ~ _T_186; // @[LZD.scala 39:27]
  assign _T_188 = _T_185 | _T_187; // @[LZD.scala 39:25]
  assign _T_189 = {_T_184,_T_188}; // @[Cat.scala 29:58]
  assign _T_190 = _T_182[1:0]; // @[LZD.scala 44:32]
  assign _T_191 = _T_190 != 2'h0; // @[LZD.scala 39:14]
  assign _T_192 = _T_190[1]; // @[LZD.scala 39:21]
  assign _T_193 = _T_190[0]; // @[LZD.scala 39:30]
  assign _T_194 = ~ _T_193; // @[LZD.scala 39:27]
  assign _T_195 = _T_192 | _T_194; // @[LZD.scala 39:25]
  assign _T_196 = {_T_191,_T_195}; // @[Cat.scala 29:58]
  assign _T_197 = _T_189[1]; // @[Shift.scala 12:21]
  assign _T_198 = _T_196[1]; // @[Shift.scala 12:21]
  assign _T_199 = _T_197 | _T_198; // @[LZD.scala 49:16]
  assign _T_200 = ~ _T_198; // @[LZD.scala 49:27]
  assign _T_201 = _T_197 | _T_200; // @[LZD.scala 49:25]
  assign _T_202 = _T_189[0:0]; // @[LZD.scala 49:47]
  assign _T_203 = _T_196[0:0]; // @[LZD.scala 49:59]
  assign _T_204 = _T_197 ? _T_202 : _T_203; // @[LZD.scala 49:35]
  assign _T_206 = {_T_199,_T_201,_T_204}; // @[Cat.scala 29:58]
  assign _T_207 = _T_181[2]; // @[Shift.scala 12:21]
  assign _T_208 = _T_206[2]; // @[Shift.scala 12:21]
  assign _T_209 = _T_207 | _T_208; // @[LZD.scala 49:16]
  assign _T_210 = ~ _T_208; // @[LZD.scala 49:27]
  assign _T_211 = _T_207 | _T_210; // @[LZD.scala 49:25]
  assign _T_212 = _T_181[1:0]; // @[LZD.scala 49:47]
  assign _T_213 = _T_206[1:0]; // @[LZD.scala 49:59]
  assign _T_214 = _T_207 ? _T_212 : _T_213; // @[LZD.scala 49:35]
  assign _T_216 = {_T_209,_T_211,_T_214}; // @[Cat.scala 29:58]
  assign _T_217 = _T_155[3:0]; // @[LZD.scala 44:32]
  assign _T_218 = _T_217[3:2]; // @[LZD.scala 43:32]
  assign _T_219 = _T_218 != 2'h0; // @[LZD.scala 39:14]
  assign _T_220 = _T_218[1]; // @[LZD.scala 39:21]
  assign _T_221 = _T_218[0]; // @[LZD.scala 39:30]
  assign _T_222 = ~ _T_221; // @[LZD.scala 39:27]
  assign _T_223 = _T_220 | _T_222; // @[LZD.scala 39:25]
  assign _T_224 = {_T_219,_T_223}; // @[Cat.scala 29:58]
  assign _T_225 = _T_217[1:0]; // @[LZD.scala 44:32]
  assign _T_226 = _T_225 != 2'h0; // @[LZD.scala 39:14]
  assign _T_227 = _T_225[1]; // @[LZD.scala 39:21]
  assign _T_228 = _T_225[0]; // @[LZD.scala 39:30]
  assign _T_229 = ~ _T_228; // @[LZD.scala 39:27]
  assign _T_230 = _T_227 | _T_229; // @[LZD.scala 39:25]
  assign _T_231 = {_T_226,_T_230}; // @[Cat.scala 29:58]
  assign _T_232 = _T_224[1]; // @[Shift.scala 12:21]
  assign _T_233 = _T_231[1]; // @[Shift.scala 12:21]
  assign _T_234 = _T_232 | _T_233; // @[LZD.scala 49:16]
  assign _T_235 = ~ _T_233; // @[LZD.scala 49:27]
  assign _T_236 = _T_232 | _T_235; // @[LZD.scala 49:25]
  assign _T_237 = _T_224[0:0]; // @[LZD.scala 49:47]
  assign _T_238 = _T_231[0:0]; // @[LZD.scala 49:59]
  assign _T_239 = _T_232 ? _T_237 : _T_238; // @[LZD.scala 49:35]
  assign _T_241 = {_T_234,_T_236,_T_239}; // @[Cat.scala 29:58]
  assign _T_242 = _T_216[3]; // @[Shift.scala 12:21]
  assign _T_244 = _T_216[2:0]; // @[LZD.scala 55:32]
  assign _T_245 = _T_242 ? _T_244 : _T_241; // @[LZD.scala 55:20]
  assign _T_246 = {_T_242,_T_245}; // @[Cat.scala 29:58]
  assign _T_247 = ~ _T_246; // @[convert.scala 21:22]
  assign _T_248 = io_B[10:0]; // @[convert.scala 22:36]
  assign _T_249 = _T_247 < 4'hb; // @[Shift.scala 16:24]
  assign _T_251 = _T_247[3]; // @[Shift.scala 12:21]
  assign _T_252 = _T_248[2:0]; // @[Shift.scala 64:52]
  assign _T_254 = {_T_252,8'h0}; // @[Cat.scala 29:58]
  assign _T_255 = _T_251 ? _T_254 : _T_248; // @[Shift.scala 64:27]
  assign _T_256 = _T_247[2:0]; // @[Shift.scala 66:70]
  assign _T_257 = _T_256[2]; // @[Shift.scala 12:21]
  assign _T_258 = _T_255[6:0]; // @[Shift.scala 64:52]
  assign _T_260 = {_T_258,4'h0}; // @[Cat.scala 29:58]
  assign _T_261 = _T_257 ? _T_260 : _T_255; // @[Shift.scala 64:27]
  assign _T_262 = _T_256[1:0]; // @[Shift.scala 66:70]
  assign _T_263 = _T_262[1]; // @[Shift.scala 12:21]
  assign _T_264 = _T_261[8:0]; // @[Shift.scala 64:52]
  assign _T_266 = {_T_264,2'h0}; // @[Cat.scala 29:58]
  assign _T_267 = _T_263 ? _T_266 : _T_261; // @[Shift.scala 64:27]
  assign _T_268 = _T_262[0:0]; // @[Shift.scala 66:70]
  assign _T_270 = _T_267[9:0]; // @[Shift.scala 64:52]
  assign _T_271 = {_T_270,1'h0}; // @[Cat.scala 29:58]
  assign _T_272 = _T_268 ? _T_271 : _T_267; // @[Shift.scala 64:27]
  assign _T_273 = _T_249 ? _T_272 : 11'h0; // @[Shift.scala 16:10]
  assign _T_274 = _T_273[10:10]; // @[convert.scala 23:34]
  assign decB_fraction = _T_273[9:0]; // @[convert.scala 24:34]
  assign _T_276 = _T_152 == 1'h0; // @[convert.scala 25:26]
  assign _T_278 = _T_152 ? _T_247 : _T_246; // @[convert.scala 25:42]
  assign _T_281 = ~ _T_274; // @[convert.scala 26:67]
  assign _T_282 = _T_150 ? _T_281 : _T_274; // @[convert.scala 26:51]
  assign _T_283 = {_T_276,_T_278,_T_282}; // @[Cat.scala 29:58]
  assign _T_285 = io_B[12:0]; // @[convert.scala 29:56]
  assign _T_286 = _T_285 != 13'h0; // @[convert.scala 29:60]
  assign _T_287 = ~ _T_286; // @[convert.scala 29:41]
  assign decB_isNaR = _T_150 & _T_287; // @[convert.scala 29:39]
  assign _T_290 = _T_150 == 1'h0; // @[convert.scala 30:19]
  assign decB_isZero = _T_290 & _T_287; // @[convert.scala 30:41]
  assign decB_scale = $signed(_T_283); // @[convert.scala 32:24]
  assign _T_299 = _T_1 ? 3'h7 : 3'h0; // @[Bitwise.scala 71:12]
  assign _T_300 = ~ _T_1; // @[PositDivisionSqrt.scala 80:40]
  assign sigA_S = {_T_299,_T_300,decA_fraction}; // @[Cat.scala 29:58]
  assign _T_302 = ~ _T_150; // @[PositDivisionSqrt.scala 82:31]
  assign sigB_S = {_T_150,_T_302,decB_fraction,2'h0}; // @[Cat.scala 29:58]
  assign _T_305 = decA_isNaR == 1'h0; // @[PositDivisionSqrt.scala 85:25]
  assign invalidSqrt = _T_305 & _T_1; // @[PositDivisionSqrt.scala 85:37]
  assign _T_306 = decA_isNaR | invalidSqrt; // @[PositDivisionSqrt.scala 88:42]
  assign _T_307 = decA_isNaR | decB_isNaR; // @[PositDivisionSqrt.scala 89:42]
  assign _T_308 = _T_307 | decB_isZero; // @[PositDivisionSqrt.scala 89:56]
  assign _T_309 = decB_isZero == 1'h0; // @[PositDivisionSqrt.scala 94:46]
  assign _T_310 = decA_isZero & _T_309; // @[PositDivisionSqrt.scala 94:43]
  assign _T_311 = decB_isNaR == 1'h0; // @[PositDivisionSqrt.scala 94:62]
  assign _T_312 = _T_310 & _T_311; // @[PositDivisionSqrt.scala 94:59]
  assign specialCaseA_S = decA_isNaR | decA_isZero; // @[PositDivisionSqrt.scala 97:38]
  assign specialCaseB_S = decB_isNaR | decB_isZero; // @[PositDivisionSqrt.scala 98:38]
  assign _T_313 = specialCaseA_S == 1'h0; // @[PositDivisionSqrt.scala 99:27]
  assign _T_314 = specialCaseB_S == 1'h0; // @[PositDivisionSqrt.scala 99:46]
  assign normalCase_S_div = _T_313 & _T_314; // @[PositDivisionSqrt.scala 99:43]
  assign normalCase_S_sqrt = _T_313 & _T_141; // @[PositDivisionSqrt.scala 100:43]
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div; // @[PositDivisionSqrt.scala 101:30]
  assign sExpQuot_S_div = $signed(decA_scale) - $signed(decB_scale); // @[PositDivisionSqrt.scala 103:38]
  assign _T_317 = decA_scale[0]; // @[PositDivisionSqrt.scala 104:50]
  assign oddSqrt_S = io_sqrtOp & _T_317; // @[PositDivisionSqrt.scala 104:37]
  assign idle = cycleNum == 4'h0; // @[PositDivisionSqrt.scala 109:39]
  assign ready = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 110:39]
  assign entering = ready & io_inValid; // @[PositDivisionSqrt.scala 111:35]
  assign entering_normalCase = entering & normalCase_S; // @[PositDivisionSqrt.scala 112:38]
  assign _T_318 = sigX_Z[13]; // @[PositDivisionSqrt.scala 113:35]
  assign _T_319 = sigX_Z[11]; // @[PositDivisionSqrt.scala 113:58]
  assign scaleNotChange = _T_318 ^ _T_319; // @[PositDivisionSqrt.scala 113:50]
  assign _T_320 = cycleNum == 4'h3; // @[PositDivisionSqrt.scala 114:39]
  assign skipCycle2 = _T_320 & scaleNotChange; // @[PositDivisionSqrt.scala 114:48]
  assign _T_321 = idle == 1'h0; // @[PositDivisionSqrt.scala 116:8]
  assign _T_322 = _T_321 | io_inValid; // @[PositDivisionSqrt.scala 116:14]
  assign _T_323 = normalCase_S == 1'h0; // @[PositDivisionSqrt.scala 117:32]
  assign _T_324 = entering & _T_323; // @[PositDivisionSqrt.scala 117:30]
  assign _T_326 = io_sqrtOp ? 4'hc : 4'he; // @[PositDivisionSqrt.scala 119:26]
  assign _T_327 = entering_normalCase ? _T_326 : 4'h0; // @[PositDivisionSqrt.scala 118:20]
  assign _GEN_9 = {{3'd0}, _T_324}; // @[PositDivisionSqrt.scala 117:64]
  assign _T_328 = _GEN_9 | _T_327; // @[PositDivisionSqrt.scala 117:64]
  assign _T_330 = skipCycle2 == 1'h0; // @[PositDivisionSqrt.scala 123:30]
  assign _T_331 = _T_321 & _T_330; // @[PositDivisionSqrt.scala 123:27]
  assign _T_333 = cycleNum - 4'h1; // @[PositDivisionSqrt.scala 123:52]
  assign _T_334 = _T_331 ? _T_333 : 4'h0; // @[PositDivisionSqrt.scala 123:20]
  assign _T_335 = _T_328 | _T_334; // @[PositDivisionSqrt.scala 122:64]
  assign _T_337 = _T_321 & skipCycle2; // @[PositDivisionSqrt.scala 124:27]
  assign _GEN_10 = {{3'd0}, _T_337}; // @[PositDivisionSqrt.scala 123:64]
  assign _T_339 = _T_335 | _GEN_10; // @[PositDivisionSqrt.scala 123:64]
  assign _T_340 = decA_scale[5:1]; // @[PositDivisionSqrt.scala 134:42]
  assign _T_342 = io_sqrtOp == 1'h0; // @[PositDivisionSqrt.scala 137:31]
  assign _T_343 = entering_normalCase & _T_342; // @[PositDivisionSqrt.scala 137:28]
  assign _T_344 = 16'h1 << cycleNum; // @[PositDivisionSqrt.scala 146:22]
  assign _T_345 = _T_344[15:2]; // @[PositDivisionSqrt.scala 146:35]
  assign _T_346 = oddSqrt_S == 1'h0; // @[PositDivisionSqrt.scala 148:26]
  assign _T_347 = ready & _T_346; // @[PositDivisionSqrt.scala 148:23]
  assign _T_348 = _T_347 ? sigA_S : 14'h0; // @[PositDivisionSqrt.scala 148:16]
  assign _T_349 = ready & oddSqrt_S; // @[PositDivisionSqrt.scala 149:23]
  assign _T_350 = {sigA_S, 1'h0}; // @[PositDivisionSqrt.scala 149:46]
  assign _T_351 = _T_350[13:0]; // @[PositDivisionSqrt.scala 149:56]
  assign _T_352 = _T_349 ? _T_351 : 14'h0; // @[PositDivisionSqrt.scala 149:16]
  assign _T_353 = _T_348 | _T_352; // @[PositDivisionSqrt.scala 148:66]
  assign _T_354 = ready == 1'h0; // @[PositDivisionSqrt.scala 150:17]
  assign _T_355 = _T_354 ? rem_Z : 14'h0; // @[PositDivisionSqrt.scala 150:16]
  assign rem = _T_353 | _T_355; // @[PositDivisionSqrt.scala 149:66]
  assign _T_357 = ready & _T_342; // @[PositDivisionSqrt.scala 152:29]
  assign _T_358 = _T_357 ? sigB_S : 14'h0; // @[PositDivisionSqrt.scala 152:22]
  assign _T_359 = ready & io_sqrtOp; // @[PositDivisionSqrt.scala 153:29]
  assign _T_360 = _T_359 ? 11'h400 : 11'h0; // @[PositDivisionSqrt.scala 153:22]
  assign _GEN_11 = {{3'd0}, _T_360}; // @[PositDivisionSqrt.scala 152:93]
  assign _T_361 = _T_358 | _GEN_11; // @[PositDivisionSqrt.scala 152:93]
  assign _T_363 = sqrtOp_Z == 1'h0; // @[PositDivisionSqrt.scala 154:33]
  assign _T_364 = _T_354 & _T_363; // @[PositDivisionSqrt.scala 154:30]
  assign _T_365 = ~ signB_Z; // @[PositDivisionSqrt.scala 154:57]
  assign _T_368 = {signB_Z,_T_365,fractB_Z,2'h0}; // @[Cat.scala 29:58]
  assign _T_369 = _T_364 ? _T_368 : 14'h0; // @[PositDivisionSqrt.scala 154:22]
  assign _T_370 = _T_361 | _T_369; // @[PositDivisionSqrt.scala 153:93]
  assign _T_372 = _T_354 & sqrtOp_Z; // @[PositDivisionSqrt.scala 155:30]
  assign _T_373 = rem[13:13]; // @[PositDivisionSqrt.scala 156:79]
  assign _T_375 = _T_373 ? 10'h3ff : 10'h0; // @[Bitwise.scala 71:12]
  assign bitMask = _T_345[12:0]; // @[PositDivisionSqrt.scala 145:21 PositDivisionSqrt.scala 146:14]
  assign _GEN_12 = {{3'd0}, _T_375}; // @[PositDivisionSqrt.scala 156:53]
  assign _T_376 = bitMask & _GEN_12; // @[PositDivisionSqrt.scala 156:53]
  assign _GEN_13 = {{1'd0}, _T_376}; // @[PositDivisionSqrt.scala 155:51]
  assign _T_377 = sigX_Z | _GEN_13; // @[PositDivisionSqrt.scala 155:51]
  assign _T_378 = bitMask[12:1]; // @[PositDivisionSqrt.scala 157:53]
  assign _GEN_14 = {{2'd0}, _T_378}; // @[PositDivisionSqrt.scala 156:85]
  assign _T_379 = _T_377 | _GEN_14; // @[PositDivisionSqrt.scala 156:85]
  assign _T_380 = _T_372 ? _T_379 : 14'h0; // @[PositDivisionSqrt.scala 155:22]
  assign trialTerm = _T_370 | _T_380; // @[PositDivisionSqrt.scala 154:93]
  assign _T_382 = trialTerm[13:13]; // @[PositDivisionSqrt.scala 162:56]
  assign _T_383 = _T_373 ^ _T_382; // @[PositDivisionSqrt.scala 162:40]
  assign _T_386 = rem + trialTerm; // @[PositDivisionSqrt.scala 163:97]
  assign _T_388 = rem - trialTerm; // @[PositDivisionSqrt.scala 164:97]
  assign _T_389 = _T_383 ? _T_386 : _T_388; // @[PositDivisionSqrt.scala 161:92]
  assign _T_394 = {rem, 1'h0}; // @[PositDivisionSqrt.scala 168:98]
  assign _T_395 = _T_394[13:0]; // @[PositDivisionSqrt.scala 168:108]
  assign _T_397 = _T_395 + trialTerm; // @[PositDivisionSqrt.scala 168:112]
  assign _T_401 = _T_395 - trialTerm; // @[PositDivisionSqrt.scala 169:112]
  assign _T_402 = _T_383 ? _T_397 : _T_401; // @[PositDivisionSqrt.scala 166:26]
  assign trialRem = ready ? _T_389 : _T_402; // @[PositDivisionSqrt.scala 159:27]
  assign _T_403 = trialRem != 14'h0; // @[PositDivisionSqrt.scala 173:35]
  assign trIsZero = _T_403 == 1'h0; // @[PositDivisionSqrt.scala 173:25]
  assign _T_404 = rem != 14'h0; // @[PositDivisionSqrt.scala 174:30]
  assign remIsZero = _T_404 == 1'h0; // @[PositDivisionSqrt.scala 174:25]
  assign _T_406 = trialRem[13:13]; // @[PositDivisionSqrt.scala 176:64]
  assign _T_407 = _T_382 ^ _T_406; // @[PositDivisionSqrt.scala 176:49]
  assign _T_408 = ~ _T_407; // @[PositDivisionSqrt.scala 176:29]
  assign _T_409 = sigX_Z[13:13]; // @[PositDivisionSqrt.scala 178:61]
  assign _T_410 = ~ _T_409; // @[PositDivisionSqrt.scala 178:49]
  assign _T_412 = remIsZero ? _T_409 : _T_408; // @[Mux.scala 87:16]
  assign newBit = trIsZero ? _T_410 : _T_412; // @[Mux.scala 87:16]
  assign _T_413 = cycleNum > 4'h2; // @[PositDivisionSqrt.scala 183:41]
  assign _T_414 = remIsZero == 1'h0; // @[PositDivisionSqrt.scala 183:51]
  assign _T_415 = _T_413 & _T_414; // @[PositDivisionSqrt.scala 183:48]
  assign _T_416 = entering_normalCase | _T_415; // @[PositDivisionSqrt.scala 183:28]
  assign _T_419 = _T_354 & newBit; // @[PositDivisionSqrt.scala 187:39]
  assign _T_420 = entering_normalCase | _T_419; // @[PositDivisionSqrt.scala 187:28]
  assign _T_423 = {newBit, 13'h0}; // @[PositDivisionSqrt.scala 188:47]
  assign _T_424 = _T_357 ? _T_423 : 14'h0; // @[PositDivisionSqrt.scala 188:18]
  assign _T_426 = _T_359 ? 12'h800 : 12'h0; // @[PositDivisionSqrt.scala 189:18]
  assign _GEN_15 = {{2'd0}, _T_426}; // @[PositDivisionSqrt.scala 188:72]
  assign _T_427 = _T_424 | _GEN_15; // @[PositDivisionSqrt.scala 188:72]
  assign _GEN_16 = {{1'd0}, bitMask}; // @[PositDivisionSqrt.scala 190:47]
  assign _T_429 = sigX_Z | _GEN_16; // @[PositDivisionSqrt.scala 190:47]
  assign _T_430 = _T_354 ? _T_429 : 14'h0; // @[PositDivisionSqrt.scala 190:18]
  assign _T_431 = _T_427 | _T_430; // @[PositDivisionSqrt.scala 189:72]
  assign _T_433 = {_T_409, 1'h0}; // @[PositDivisionSqrt.scala 196:53]
  assign sigXBias = scaleNotChange ? _T_433 : {{1'd0}, _T_409}; // @[PositDivisionSqrt.scala 196:21]
  assign _GEN_17 = {{12'd0}, sigXBias}; // @[PositDivisionSqrt.scala 197:25]
  assign realSigX = sigX_Z + _GEN_17; // @[PositDivisionSqrt.scala 197:25]
  assign _T_436 = realSigX[10:1]; // @[PositDivisionSqrt.scala 200:97]
  assign _T_437 = realSigX[9:0]; // @[PositDivisionSqrt.scala 201:97]
  assign realFrac = scaleNotChange ? _T_436 : _T_437; // @[PositDivisionSqrt.scala 198:21]
  assign _T_438 = realSigX[13]; // @[PositDivisionSqrt.scala 205:33]
  assign _T_439 = realSigX[11]; // @[PositDivisionSqrt.scala 205:58]
  assign _T_440 = _T_438 ^ _T_439; // @[PositDivisionSqrt.scala 205:48]
  assign scaleNeedSub = ~ _T_440; // @[PositDivisionSqrt.scala 205:23]
  assign _T_442 = realSigX[10]; // @[PositDivisionSqrt.scala 206:56]
  assign notNeedSubTwo = _T_438 ^ _T_442; // @[PositDivisionSqrt.scala 206:46]
  assign scaleSubOne = scaleNeedSub & notNeedSubTwo; // @[PositDivisionSqrt.scala 207:36]
  assign _T_443 = ~ notNeedSubTwo; // @[PositDivisionSqrt.scala 208:38]
  assign scaleSubTwo = scaleNeedSub & _T_443; // @[PositDivisionSqrt.scala 208:36]
  assign _T_444 = {scaleSubTwo,scaleSubOne}; // @[Cat.scala 29:58]
  assign _T_445 = {1'b0,$signed(_T_444)}; // @[PositDivisionSqrt.scala 209:63]
  assign _GEN_18 = {{4{_T_445[2]}},_T_445}; // @[PositDivisionSqrt.scala 209:31]
  assign _T_447 = $signed(scale_Z) - $signed(_GEN_18); // @[PositDivisionSqrt.scala 209:31]
  assign realExp = $signed(_T_447); // @[PositDivisionSqrt.scala 209:31]
  assign underflow = $signed(realExp) < $signed(-7'sh18); // @[PositDivisionSqrt.scala 210:31]
  assign overflow = $signed(realExp) > $signed(7'sh18); // @[PositDivisionSqrt.scala 211:31]
  assign decQ_sign = realSigX[13:13]; // @[PositDivisionSqrt.scala 215:33]
  assign _T_449 = underflow ? $signed(-7'sh18) : $signed(realExp); // @[Mux.scala 87:16]
  assign _T_450 = overflow ? $signed(7'sh18) : $signed(_T_449); // @[Mux.scala 87:16]
  assign outValid = cycleNum == 4'h1; // @[PositDivisionSqrt.scala 229:28]
  assign _GEN_19 = _T_450[5:0]; // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign decQ_scale = $signed(_GEN_19); // @[PositDivisionSqrt.scala 204:27 PositDivisionSqrt.scala 216:23]
  assign _T_455 = decQ_scale[0]; // @[convert.scala 46:61]
  assign _T_456 = ~ _T_455; // @[convert.scala 46:52]
  assign _T_458 = decQ_sign ? _T_456 : _T_455; // @[convert.scala 46:42]
  assign _T_459 = decQ_scale[5:1]; // @[convert.scala 48:34]
  assign _T_460 = _T_459[4:4]; // @[convert.scala 49:36]
  assign _T_462 = ~ _T_459; // @[convert.scala 50:36]
  assign _T_463 = $signed(_T_462); // @[convert.scala 50:36]
  assign _T_464 = _T_460 ? $signed(_T_463) : $signed(_T_459); // @[convert.scala 50:28]
  assign _T_465 = _T_460 ^ decQ_sign; // @[convert.scala 51:31]
  assign _T_466 = ~ _T_465; // @[convert.scala 52:43]
  assign _T_470 = {_T_466,_T_465,_T_458,realFrac,3'h0}; // @[Cat.scala 29:58]
  assign _T_471 = $unsigned(_T_464); // @[Shift.scala 39:17]
  assign _T_472 = _T_471 < 5'h10; // @[Shift.scala 39:24]
  assign _T_473 = _T_464[3:0]; // @[Shift.scala 40:44]
  assign _T_474 = _T_470[15:8]; // @[Shift.scala 90:30]
  assign _T_475 = _T_470[7:0]; // @[Shift.scala 90:48]
  assign _T_476 = _T_475 != 8'h0; // @[Shift.scala 90:57]
  assign _GEN_20 = {{7'd0}, _T_476}; // @[Shift.scala 90:39]
  assign _T_477 = _T_474 | _GEN_20; // @[Shift.scala 90:39]
  assign _T_478 = _T_473[3]; // @[Shift.scala 12:21]
  assign _T_479 = _T_470[15]; // @[Shift.scala 12:21]
  assign _T_481 = _T_479 ? 8'hff : 8'h0; // @[Bitwise.scala 71:12]
  assign _T_482 = {_T_481,_T_477}; // @[Cat.scala 29:58]
  assign _T_483 = _T_478 ? _T_482 : _T_470; // @[Shift.scala 91:22]
  assign _T_484 = _T_473[2:0]; // @[Shift.scala 92:77]
  assign _T_485 = _T_483[15:4]; // @[Shift.scala 90:30]
  assign _T_486 = _T_483[3:0]; // @[Shift.scala 90:48]
  assign _T_487 = _T_486 != 4'h0; // @[Shift.scala 90:57]
  assign _GEN_21 = {{11'd0}, _T_487}; // @[Shift.scala 90:39]
  assign _T_488 = _T_485 | _GEN_21; // @[Shift.scala 90:39]
  assign _T_489 = _T_484[2]; // @[Shift.scala 12:21]
  assign _T_490 = _T_483[15]; // @[Shift.scala 12:21]
  assign _T_492 = _T_490 ? 4'hf : 4'h0; // @[Bitwise.scala 71:12]
  assign _T_493 = {_T_492,_T_488}; // @[Cat.scala 29:58]
  assign _T_494 = _T_489 ? _T_493 : _T_483; // @[Shift.scala 91:22]
  assign _T_495 = _T_484[1:0]; // @[Shift.scala 92:77]
  assign _T_496 = _T_494[15:2]; // @[Shift.scala 90:30]
  assign _T_497 = _T_494[1:0]; // @[Shift.scala 90:48]
  assign _T_498 = _T_497 != 2'h0; // @[Shift.scala 90:57]
  assign _GEN_22 = {{13'd0}, _T_498}; // @[Shift.scala 90:39]
  assign _T_499 = _T_496 | _GEN_22; // @[Shift.scala 90:39]
  assign _T_500 = _T_495[1]; // @[Shift.scala 12:21]
  assign _T_501 = _T_494[15]; // @[Shift.scala 12:21]
  assign _T_503 = _T_501 ? 2'h3 : 2'h0; // @[Bitwise.scala 71:12]
  assign _T_504 = {_T_503,_T_499}; // @[Cat.scala 29:58]
  assign _T_505 = _T_500 ? _T_504 : _T_494; // @[Shift.scala 91:22]
  assign _T_506 = _T_495[0:0]; // @[Shift.scala 92:77]
  assign _T_507 = _T_505[15:1]; // @[Shift.scala 90:30]
  assign _T_508 = _T_505[0:0]; // @[Shift.scala 90:48]
  assign _GEN_23 = {{14'd0}, _T_508}; // @[Shift.scala 90:39]
  assign _T_510 = _T_507 | _GEN_23; // @[Shift.scala 90:39]
  assign _T_512 = _T_505[15]; // @[Shift.scala 12:21]
  assign _T_513 = {_T_512,_T_510}; // @[Cat.scala 29:58]
  assign _T_514 = _T_506 ? _T_513 : _T_505; // @[Shift.scala 91:22]
  assign _T_517 = _T_479 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_518 = _T_472 ? _T_514 : _T_517; // @[Shift.scala 39:10]
  assign _T_519 = _T_518[3]; // @[convert.scala 55:31]
  assign _T_520 = _T_518[2]; // @[convert.scala 56:31]
  assign _T_521 = _T_518[1]; // @[convert.scala 57:31]
  assign _T_522 = _T_518[0]; // @[convert.scala 58:31]
  assign _T_523 = _T_518[15:3]; // @[convert.scala 59:69]
  assign _T_524 = _T_523 != 13'h0; // @[convert.scala 59:81]
  assign _T_525 = ~ _T_524; // @[convert.scala 59:50]
  assign _T_527 = _T_523 == 13'h1fff; // @[convert.scala 60:81]
  assign _T_528 = _T_519 | _T_521; // @[convert.scala 61:44]
  assign _T_529 = _T_528 | _T_522; // @[convert.scala 61:52]
  assign _T_530 = _T_520 & _T_529; // @[convert.scala 61:36]
  assign _T_531 = ~ _T_527; // @[convert.scala 62:63]
  assign _T_532 = _T_531 & _T_530; // @[convert.scala 62:103]
  assign _T_533 = _T_525 | _T_532; // @[convert.scala 62:60]
  assign _GEN_24 = {{12'd0}, _T_533}; // @[convert.scala 63:56]
  assign _T_536 = _T_523 + _GEN_24; // @[convert.scala 63:56]
  assign _T_537 = {decQ_sign,_T_536}; // @[Cat.scala 29:58]
  assign _T_539 = isZero_Z ? 14'h0 : _T_537; // @[Mux.scala 87:16]
  assign io_inReady = cycleNum <= 4'h1; // @[PositDivisionSqrt.scala 231:17]
  assign io_diviValid = outValid & _T_363; // @[PositDivisionSqrt.scala 232:17]
  assign io_sqrtValid = outValid & sqrtOp_Z; // @[PositDivisionSqrt.scala 233:17]
  assign io_invalidExc = isNaR_Z; // @[PositDivisionSqrt.scala 234:17]
  assign io_Q = isNaR_Z ? 14'h2000 : _T_539; // @[PositDivisionSqrt.scala 235:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sqrtOp_Z = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  isNaR_Z = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isZero_Z = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  scale_Z = _RAND_4[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  signB_Z = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fractB_Z = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rem_Z = _RAND_7[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  sigX_Z = _RAND_8[13:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      cycleNum <= 4'h0;
    end else begin
      if (_T_322) begin
        cycleNum <= _T_339;
      end
    end
    if (entering) begin
      sqrtOp_Z <= io_sqrtOp;
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isNaR_Z <= _T_306;
      end else begin
        isNaR_Z <= _T_308;
      end
    end
    if (entering) begin
      if (io_sqrtOp) begin
        isZero_Z <= decA_isZero;
      end else begin
        isZero_Z <= _T_312;
      end
    end
    if (entering_normalCase) begin
      if (io_sqrtOp) begin
        scale_Z <= {{2{_T_340[4]}},_T_340};
      end else begin
        scale_Z <= sExpQuot_S_div;
      end
    end
    if (_T_343) begin
      signB_Z <= _T_150;
    end
    if (_T_343) begin
      fractB_Z <= decB_fraction;
    end
    if (_T_416) begin
      if (ready) begin
        if (_T_383) begin
          rem_Z <= _T_386;
        end else begin
          rem_Z <= _T_388;
        end
      end else begin
        if (_T_383) begin
          rem_Z <= _T_397;
        end else begin
          rem_Z <= _T_401;
        end
      end
    end
    if (_T_420) begin
      sigX_Z <= _T_431;
    end
  end
endmodule
